// Example code for an AHBLite System-on-Chip
//  Iain McNally
//  ECS, University of Soutampton
//
// This module is an AHB-Lite Slave containing a ROM
//
// Number of addressable locations : 2**MEMWIDTH
// Size of each addressable location : 8 bits
// Supported transfer sizes : Word, Halfword, Byte
// Alignment of base address : Word aligned
//

`ifdef PROG_FILE_VMEM
  // already defined - do nothing
`else
  `define PROG_FILE_VMEM  "code.vmem"
`endif

module ahb_rom #(
  parameter MEMWIDTH = 14
)(
  //AHBLITE INTERFACE

    //Slave Select Signal
    input HSEL,
    //Global Signals
    input HCLK,
    input HRESETn,
    //Address, Control & Write Data
    input HREADY,
    input [31:0] HADDR,
    input [1:0] HTRANS,
    input HWRITE,
    input [2:0] HSIZE,
    input [31:0] HWDATA,
    // Transfer Response & Read Data
    output HREADYOUT,
    output [31:0] HRDATA

);

timeunit 1ns;
timeprecision 100ps;

  localparam No_Transfer = 2'b0;

// Memory Array  
  logic [31:0] memory[0:2293];

//control signals are stored in registers
  logic read_enable;
  logic [MEMWIDTH-3:0] word_address;
  logic [3:0] byte_select;
  

// BEGIN CUSTOM

  assign memory[ 0 ] = 32'h2000032C;
  assign memory[ 1 ] = 32'h000000C1;
  assign memory[ 2 ] = 32'h00000121;
  assign memory[ 3 ] = 32'h00000125;
  assign memory[ 4 ] = 32'h00000129;
  assign memory[ 5 ] = 32'h0000012D;
  assign memory[ 6 ] = 32'h00000131;
  assign memory[ 7 ] = 32'h00000000;
  assign memory[ 8 ] = 32'h00000000;
  assign memory[ 9 ] = 32'h00000000;
  assign memory[ 10 ] = 32'h00000000;
  assign memory[ 11 ] = 32'h00000135;
  assign memory[ 12 ] = 32'h00000139;
  assign memory[ 13 ] = 32'h00000000;
  assign memory[ 14 ] = 32'h0000013D;
  assign memory[ 15 ] = 32'h000004C9;
  assign memory[ 16 ] = 32'h00000145;
  assign memory[ 17 ] = 32'h00000145;
  assign memory[ 18 ] = 32'h00000145;
  assign memory[ 19 ] = 32'h00000145;
  assign memory[ 20 ] = 32'h00000145;
  assign memory[ 21 ] = 32'h00000145;
  assign memory[ 22 ] = 32'h00000145;
  assign memory[ 23 ] = 32'h00000145;
  assign memory[ 24 ] = 32'h00000145;
  assign memory[ 25 ] = 32'h00000145;
  assign memory[ 26 ] = 32'h00000145;
  assign memory[ 27 ] = 32'h00000145;
  assign memory[ 28 ] = 32'h00000145;
  assign memory[ 29 ] = 32'h00000149;
  assign memory[ 30 ] = 32'h0000014D;
  assign memory[ 31 ] = 32'h00000151;
  assign memory[ 32 ] = 32'h00000155;
  assign memory[ 33 ] = 32'h00000159;
  assign memory[ 34 ] = 32'h0000015D;
  assign memory[ 35 ] = 32'h00000161;
  assign memory[ 36 ] = 32'h00000165;
  assign memory[ 37 ] = 32'h00000169;
  assign memory[ 38 ] = 32'h00000000;
  assign memory[ 39 ] = 32'h00000000;
  assign memory[ 40 ] = 32'h0000016D;
  assign memory[ 41 ] = 32'h00000171;
  assign memory[ 42 ] = 32'h00000175;
  assign memory[ 43 ] = 32'h00000000;
  assign memory[ 44 ] = 32'h00000179;
  assign memory[ 45 ] = 32'h0000017D;
  assign memory[ 46 ] = 32'h00000181;
  assign memory[ 47 ] = 32'h00000185;
  assign memory[ 48 ] = 32'hB083B500;
  assign memory[ 49 ] = 32'h93004B11;
  assign memory[ 50 ] = 32'h93014B11;
  assign memory[ 51 ] = 32'h9B019A00;
  assign memory[ 52 ] = 32'hD00C429A;
  assign memory[ 53 ] = 32'h9B01E007;
  assign memory[ 54 ] = 32'h92011D1A;
  assign memory[ 55 ] = 32'h1D119A00;
  assign memory[ 56 ] = 32'h68129100;
  assign memory[ 57 ] = 32'h9A01601A;
  assign memory[ 58 ] = 32'h429A4B0A;
  assign memory[ 59 ] = 32'h4B0AD3F3;
  assign memory[ 60 ] = 32'hE0049301;
  assign memory[ 61 ] = 32'h1D1A9B01;
  assign memory[ 62 ] = 32'h22009201;
  assign memory[ 63 ] = 32'h9A01601A;
  assign memory[ 64 ] = 32'h429A4B06;
  assign memory[ 65 ] = 32'hF001D3F6;
  assign memory[ 66 ] = 32'hE7FEFC27;
  assign memory[ 67 ] = 32'h00002318;
  assign memory[ 68 ] = 32'h20000000;
  assign memory[ 69 ] = 32'h200000C0;
  assign memory[ 70 ] = 32'h200000C0;
  assign memory[ 71 ] = 32'h20000100;
  assign memory[ 72 ] = 32'h46C0E7FE;
  assign memory[ 73 ] = 32'h46C0E7FE;
  assign memory[ 74 ] = 32'h46C0E7FE;
  assign memory[ 75 ] = 32'h46C0E7FE;
  assign memory[ 76 ] = 32'h46C0E7FE;
  assign memory[ 77 ] = 32'h46C0E7FE;
  assign memory[ 78 ] = 32'h46C0E7FE;
  assign memory[ 79 ] = 32'h46C0E7FE;
  assign memory[ 80 ] = 32'h46C0E7FE;
  assign memory[ 81 ] = 32'h46C0E7FE;
  assign memory[ 82 ] = 32'h46C0E7FE;
  assign memory[ 83 ] = 32'h46C0E7FE;
  assign memory[ 84 ] = 32'h46C0E7FE;
  assign memory[ 85 ] = 32'h46C0E7FE;
  assign memory[ 86 ] = 32'h46C0E7FE;
  assign memory[ 87 ] = 32'h46C0E7FE;
  assign memory[ 88 ] = 32'h46C0E7FE;
  assign memory[ 89 ] = 32'h46C0E7FE;
  assign memory[ 90 ] = 32'h46C0E7FE;
  assign memory[ 91 ] = 32'h46C0E7FE;
  assign memory[ 92 ] = 32'h46C0E7FE;
  assign memory[ 93 ] = 32'h46C0E7FE;
  assign memory[ 94 ] = 32'h46C0E7FE;
  assign memory[ 95 ] = 32'h46C0E7FE;
  assign memory[ 96 ] = 32'h46C0E7FE;
  assign memory[ 97 ] = 32'h46C0E7FE;
  assign memory[ 98 ] = 32'h9001B082;
  assign memory[ 99 ] = 32'h9A019100;
  assign memory[ 100 ] = 32'h18D39B00;
  assign memory[ 101 ] = 32'hB0020018;
  assign memory[ 102 ] = 32'h46C04770;
  assign memory[ 103 ] = 32'h9001B082;
  assign memory[ 104 ] = 32'h9A019100;
  assign memory[ 105 ] = 32'h1AD39B00;
  assign memory[ 106 ] = 32'hB0020018;
  assign memory[ 107 ] = 32'h46C04770;
  assign memory[ 108 ] = 32'hB083B5F0;
  assign memory[ 109 ] = 32'h91009001;
  assign memory[ 110 ] = 32'h000A9901;
  assign memory[ 111 ] = 32'h000B17C9;
  assign memory[ 112 ] = 32'h039D0C91;
  assign memory[ 113 ] = 32'h0394430D;
  assign memory[ 114 ] = 32'h001E9B00;
  assign memory[ 115 ] = 32'h001F17DB;
  assign memory[ 116 ] = 32'h003B0032;
  assign memory[ 117 ] = 32'h00290020;
  assign memory[ 118 ] = 32'hFEC4F001;
  assign memory[ 119 ] = 32'h000C0003;
  assign memory[ 120 ] = 32'hB0030018;
  assign memory[ 121 ] = 32'h46C0BDF0;
  assign memory[ 122 ] = 32'h681B4B04;
  assign memory[ 123 ] = 32'h681B3304;
  assign memory[ 124 ] = 32'h41931E5A;
  assign memory[ 125 ] = 32'h0018B2DB;
  assign memory[ 126 ] = 32'h46C04770;
  assign memory[ 127 ] = 32'h20000000;
  assign memory[ 128 ] = 32'h681B4B02;
  assign memory[ 129 ] = 32'h0018681B;
  assign memory[ 130 ] = 32'h46C04770;
  assign memory[ 131 ] = 32'h20000000;
  assign memory[ 132 ] = 32'h4B0446C0;
  assign memory[ 133 ] = 32'h3304681B;
  assign memory[ 134 ] = 32'h2B00681B;
  assign memory[ 135 ] = 32'h46C0D0F9;
  assign memory[ 136 ] = 32'h46C04770;
  assign memory[ 137 ] = 32'h20000000;
  assign memory[ 138 ] = 32'h681B4B05;
  assign memory[ 139 ] = 32'h681B3318;
  assign memory[ 140 ] = 32'h40132201;
  assign memory[ 141 ] = 32'h41931E5A;
  assign memory[ 142 ] = 32'h0018B2DB;
  assign memory[ 143 ] = 32'h46C04770;
  assign memory[ 144 ] = 32'h20000008;
  assign memory[ 145 ] = 32'h681B4B05;
  assign memory[ 146 ] = 32'h681B3318;
  assign memory[ 147 ] = 32'h40132202;
  assign memory[ 148 ] = 32'h41931E5A;
  assign memory[ 149 ] = 32'h0018B2DB;
  assign memory[ 150 ] = 32'h46C04770;
  assign memory[ 151 ] = 32'h20000008;
  assign memory[ 152 ] = 32'h9001B082;
  assign memory[ 153 ] = 32'h681B4B03;
  assign memory[ 154 ] = 32'h601A9A01;
  assign memory[ 155 ] = 32'hB00246C0;
  assign memory[ 156 ] = 32'h46C04770;
  assign memory[ 157 ] = 32'h20000008;
  assign memory[ 158 ] = 32'h681B4B02;
  assign memory[ 159 ] = 32'h0018681B;
  assign memory[ 160 ] = 32'h46C04770;
  assign memory[ 161 ] = 32'h20000008;
  assign memory[ 162 ] = 32'hB085B530;
  assign memory[ 163 ] = 32'h000C0005;
  assign memory[ 164 ] = 32'h00190010;
  assign memory[ 165 ] = 32'h3307466B;
  assign memory[ 166 ] = 32'h701A1C2A;
  assign memory[ 167 ] = 32'h3306466B;
  assign memory[ 168 ] = 32'h701A1C22;
  assign memory[ 169 ] = 32'h3305466B;
  assign memory[ 170 ] = 32'h701A1C02;
  assign memory[ 171 ] = 32'h1C0AAB01;
  assign memory[ 172 ] = 32'h2300701A;
  assign memory[ 173 ] = 32'h466B9303;
  assign memory[ 174 ] = 32'h781B3307;
  assign memory[ 175 ] = 32'h466B061A;
  assign memory[ 176 ] = 32'h781B3306;
  assign memory[ 177 ] = 32'h18D2041B;
  assign memory[ 178 ] = 32'h3305466B;
  assign memory[ 179 ] = 32'h021B781B;
  assign memory[ 180 ] = 32'hAB0118D2;
  assign memory[ 181 ] = 32'h18D3781B;
  assign memory[ 182 ] = 32'h4B049303;
  assign memory[ 183 ] = 32'h3304681B;
  assign memory[ 184 ] = 32'h601A9A03;
  assign memory[ 185 ] = 32'hB00546C0;
  assign memory[ 186 ] = 32'h46C0BD30;
  assign memory[ 187 ] = 32'h20000008;
  assign memory[ 188 ] = 32'h681B4B02;
  assign memory[ 189 ] = 32'h681B3304;
  assign memory[ 190 ] = 32'h47700018;
  assign memory[ 191 ] = 32'h20000008;
  assign memory[ 192 ] = 32'h681B4B02;
  assign memory[ 193 ] = 32'h681B3308;
  assign memory[ 194 ] = 32'h47700018;
  assign memory[ 195 ] = 32'h20000008;
  assign memory[ 196 ] = 32'h681B4B02;
  assign memory[ 197 ] = 32'h681B330C;
  assign memory[ 198 ] = 32'h47700018;
  assign memory[ 199 ] = 32'h20000008;
  assign memory[ 200 ] = 32'h681B4B02;
  assign memory[ 201 ] = 32'h681B3310;
  assign memory[ 202 ] = 32'h47700018;
  assign memory[ 203 ] = 32'h20000008;
  assign memory[ 204 ] = 32'hB085B530;
  assign memory[ 205 ] = 32'h000C0005;
  assign memory[ 206 ] = 32'h00190010;
  assign memory[ 207 ] = 32'h3307466B;
  assign memory[ 208 ] = 32'h701A1C2A;
  assign memory[ 209 ] = 32'h3306466B;
  assign memory[ 210 ] = 32'h701A1C22;
  assign memory[ 211 ] = 32'h3305466B;
  assign memory[ 212 ] = 32'h701A1C02;
  assign memory[ 213 ] = 32'h1C0AAB01;
  assign memory[ 214 ] = 32'h2300701A;
  assign memory[ 215 ] = 32'h466B9303;
  assign memory[ 216 ] = 32'h781B3307;
  assign memory[ 217 ] = 32'h466B061A;
  assign memory[ 218 ] = 32'h781B3306;
  assign memory[ 219 ] = 32'h18D2041B;
  assign memory[ 220 ] = 32'h3305466B;
  assign memory[ 221 ] = 32'h021B781B;
  assign memory[ 222 ] = 32'hAB0118D2;
  assign memory[ 223 ] = 32'h18D3781B;
  assign memory[ 224 ] = 32'h4B049303;
  assign memory[ 225 ] = 32'h3310681B;
  assign memory[ 226 ] = 32'h601A9A03;
  assign memory[ 227 ] = 32'hB00546C0;
  assign memory[ 228 ] = 32'h46C0BD30;
  assign memory[ 229 ] = 32'h20000008;
  assign memory[ 230 ] = 32'h9001B084;
  assign memory[ 231 ] = 32'h23009100;
  assign memory[ 232 ] = 32'h9B019303;
  assign memory[ 233 ] = 32'h9B039303;
  assign memory[ 234 ] = 32'h93033302;
  assign memory[ 235 ] = 32'h009B9B00;
  assign memory[ 236 ] = 32'h18D39A03;
  assign memory[ 237 ] = 32'h4B049303;
  assign memory[ 238 ] = 32'h3314681B;
  assign memory[ 239 ] = 32'h601A9A03;
  assign memory[ 240 ] = 32'hB00446C0;
  assign memory[ 241 ] = 32'h46C04770;
  assign memory[ 242 ] = 32'h20000008;
  assign memory[ 243 ] = 32'h9001B082;
  assign memory[ 244 ] = 32'h681B4B03;
  assign memory[ 245 ] = 32'h601A9A01;
  assign memory[ 246 ] = 32'hB00246C0;
  assign memory[ 247 ] = 32'h46C04770;
  assign memory[ 248 ] = 32'h20000004;
  assign memory[ 249 ] = 32'h9001B082;
  assign memory[ 250 ] = 32'h681B4B03;
  assign memory[ 251 ] = 32'h9A013304;
  assign memory[ 252 ] = 32'h46C0601A;
  assign memory[ 253 ] = 32'h4770B002;
  assign memory[ 254 ] = 32'h20000004;
  assign memory[ 255 ] = 32'h681B4B02;
  assign memory[ 256 ] = 32'h0018681B;
  assign memory[ 257 ] = 32'h46C04770;
  assign memory[ 258 ] = 32'h20000004;
  assign memory[ 259 ] = 32'h681B4B02;
  assign memory[ 260 ] = 32'h681B3304;
  assign memory[ 261 ] = 32'h47700018;
  assign memory[ 262 ] = 32'h20000004;
  assign memory[ 263 ] = 32'hB084B510;
  assign memory[ 264 ] = 32'h00080004;
  assign memory[ 265 ] = 32'h466B0011;
  assign memory[ 266 ] = 32'h1C223307;
  assign memory[ 267 ] = 32'h466B701A;
  assign memory[ 268 ] = 32'h1C023306;
  assign memory[ 269 ] = 32'h466B701A;
  assign memory[ 270 ] = 32'h1C0A3305;
  assign memory[ 271 ] = 32'h466B701A;
  assign memory[ 272 ] = 32'h781B3307;
  assign memory[ 273 ] = 32'h466B025A;
  assign memory[ 274 ] = 32'h781B3306;
  assign memory[ 275 ] = 32'h18D2021B;
  assign memory[ 276 ] = 32'h3305466B;
  assign memory[ 277 ] = 32'h18D3781B;
  assign memory[ 278 ] = 32'h4B049303;
  assign memory[ 279 ] = 32'h3308681B;
  assign memory[ 280 ] = 32'h601A9A03;
  assign memory[ 281 ] = 32'hB00446C0;
  assign memory[ 282 ] = 32'h46C0BD10;
  assign memory[ 283 ] = 32'h20000004;
  assign memory[ 284 ] = 32'h681B4B02;
  assign memory[ 285 ] = 32'h681B3308;
  assign memory[ 286 ] = 32'h47700018;
  assign memory[ 287 ] = 32'h20000004;
  assign memory[ 288 ] = 32'h0002B084;
  assign memory[ 289 ] = 32'h3307466B;
  assign memory[ 290 ] = 32'h2300701A;
  assign memory[ 291 ] = 32'h466B9303;
  assign memory[ 292 ] = 32'h781B3307;
  assign memory[ 293 ] = 32'h9B039303;
  assign memory[ 294 ] = 32'h93033302;
  assign memory[ 295 ] = 32'h681B4B03;
  assign memory[ 296 ] = 32'h9A03330C;
  assign memory[ 297 ] = 32'h46C0601A;
  assign memory[ 298 ] = 32'h4770B004;
  assign memory[ 299 ] = 32'h20000004;
  assign memory[ 300 ] = 32'h681B4B04;
  assign memory[ 301 ] = 32'h681B3310;
  assign memory[ 302 ] = 32'h41931E5A;
  assign memory[ 303 ] = 32'h0018B2DB;
  assign memory[ 304 ] = 32'h46C04770;
  assign memory[ 305 ] = 32'h20000004;
  assign memory[ 306 ] = 32'h681B4B03;
  assign memory[ 307 ] = 32'h4B021C5A;
  assign memory[ 308 ] = 32'h46C0601A;
  assign memory[ 309 ] = 32'h46C04770;
  assign memory[ 310 ] = 32'h200000C0;
  assign memory[ 311 ] = 32'h9001B082;
  assign memory[ 312 ] = 32'h9A014B06;
  assign memory[ 313 ] = 32'h605A3A01;
  assign memory[ 314 ] = 32'h22004B04;
  assign memory[ 315 ] = 32'h4B03609A;
  assign memory[ 316 ] = 32'h601A2207;
  assign memory[ 317 ] = 32'hB00246C0;
  assign memory[ 318 ] = 32'h46C04770;
  assign memory[ 319 ] = 32'hE000E010;
  assign memory[ 320 ] = 32'h9001B084;
  assign memory[ 321 ] = 32'h681B4B06;
  assign memory[ 322 ] = 32'h9B019303;
  assign memory[ 323 ] = 32'hD0022B00;
  assign memory[ 324 ] = 32'h9A039B01;
  assign memory[ 325 ] = 32'h9B03601A;
  assign memory[ 326 ] = 32'hB0040018;
  assign memory[ 327 ] = 32'h46C04770;
  assign memory[ 328 ] = 32'h200000C0;
  assign memory[ 329 ] = 32'hB085B500;
  assign memory[ 330 ] = 32'h4B119001;
  assign memory[ 331 ] = 32'h9303689B;
  assign memory[ 332 ] = 32'h03DA9B01;
  assign memory[ 333 ] = 32'h009923FA;
  assign memory[ 334 ] = 32'hF0010010;
  assign memory[ 335 ] = 32'h0003FB9D;
  assign memory[ 336 ] = 32'h46C09302;
  assign memory[ 337 ] = 32'h685A4B0A;
  assign memory[ 338 ] = 32'h18D29B03;
  assign memory[ 339 ] = 32'h689B4B08;
  assign memory[ 340 ] = 32'h4B071AD2;
  assign memory[ 341 ] = 32'h0019685B;
  assign memory[ 342 ] = 32'hF0010010;
  assign memory[ 343 ] = 32'h000BFC13;
  assign memory[ 344 ] = 32'h9B02001A;
  assign memory[ 345 ] = 32'hD3ED429A;
  assign memory[ 346 ] = 32'hB00546C0;
  assign memory[ 347 ] = 32'h46C0BD00;
  assign memory[ 348 ] = 32'hE000E010;
  assign memory[ 349 ] = 32'h46C0B510;
  assign memory[ 350 ] = 32'hFF9AF7FF;
  assign memory[ 351 ] = 32'hD1FB1E03;
  assign memory[ 352 ] = 32'hBD1046C0;
  assign memory[ 353 ] = 32'hB082B510;
  assign memory[ 354 ] = 32'h00080004;
  assign memory[ 355 ] = 32'h466B0011;
  assign memory[ 356 ] = 32'h1C223307;
  assign memory[ 357 ] = 32'h466B701A;
  assign memory[ 358 ] = 32'h1C023306;
  assign memory[ 359 ] = 32'h466B701A;
  assign memory[ 360 ] = 32'h1C0A3305;
  assign memory[ 361 ] = 32'hF7FF701A;
  assign memory[ 362 ] = 32'h466BFFE5;
  assign memory[ 363 ] = 32'h781A3305;
  assign memory[ 364 ] = 32'h3306466B;
  assign memory[ 365 ] = 32'h466B7819;
  assign memory[ 366 ] = 32'h781B3307;
  assign memory[ 367 ] = 32'hF7FF0018;
  assign memory[ 368 ] = 32'h2000FF2D;
  assign memory[ 369 ] = 32'hFF5CF7FF;
  assign memory[ 370 ] = 32'hB00246C0;
  assign memory[ 371 ] = 32'h46C0BD10;
  assign memory[ 372 ] = 32'hF7FFB510;
  assign memory[ 373 ] = 32'h2001FFCF;
  assign memory[ 374 ] = 32'hFF52F7FF;
  assign memory[ 375 ] = 32'hBD1046C0;
  assign memory[ 376 ] = 32'h2032B510;
  assign memory[ 377 ] = 32'hFF9EF7FF;
  assign memory[ 378 ] = 32'h21002230;
  assign memory[ 379 ] = 32'hF7FF2000;
  assign memory[ 380 ] = 32'h2000FF15;
  assign memory[ 381 ] = 32'hFF44F7FF;
  assign memory[ 382 ] = 32'hF7FF2005;
  assign memory[ 383 ] = 32'h2230FF93;
  assign memory[ 384 ] = 32'h20002100;
  assign memory[ 385 ] = 32'hFF0AF7FF;
  assign memory[ 386 ] = 32'hF7FF2000;
  assign memory[ 387 ] = 32'h2001FF39;
  assign memory[ 388 ] = 32'hFF88F7FF;
  assign memory[ 389 ] = 32'h21002230;
  assign memory[ 390 ] = 32'hF7FF2000;
  assign memory[ 391 ] = 32'h2000FEFF;
  assign memory[ 392 ] = 32'hFF2EF7FF;
  assign memory[ 393 ] = 32'hF7FF2001;
  assign memory[ 394 ] = 32'h2238FF7D;
  assign memory[ 395 ] = 32'h20002100;
  assign memory[ 396 ] = 32'hFFA8F7FF;
  assign memory[ 397 ] = 32'h21002208;
  assign memory[ 398 ] = 32'hF7FF2000;
  assign memory[ 399 ] = 32'h2201FFA3;
  assign memory[ 400 ] = 32'h20002100;
  assign memory[ 401 ] = 32'hFF9EF7FF;
  assign memory[ 402 ] = 32'h21002206;
  assign memory[ 403 ] = 32'hF7FF2000;
  assign memory[ 404 ] = 32'h220CFF99;
  assign memory[ 405 ] = 32'h20002100;
  assign memory[ 406 ] = 32'hFF94F7FF;
  assign memory[ 407 ] = 32'hBD1046C0;
  assign memory[ 408 ] = 32'h9001B084;
  assign memory[ 409 ] = 32'h2B0F9B01;
  assign memory[ 410 ] = 32'h9B01D855;
  assign memory[ 411 ] = 32'h4B2F009A;
  assign memory[ 412 ] = 32'h681B18D3;
  assign memory[ 413 ] = 32'h230F469F;
  assign memory[ 414 ] = 32'h2230446B;
  assign memory[ 415 ] = 32'hE04F701A;
  assign memory[ 416 ] = 32'h446B230F;
  assign memory[ 417 ] = 32'h701A2231;
  assign memory[ 418 ] = 32'h230FE04A;
  assign memory[ 419 ] = 32'h2232446B;
  assign memory[ 420 ] = 32'hE045701A;
  assign memory[ 421 ] = 32'h446B230F;
  assign memory[ 422 ] = 32'h701A2233;
  assign memory[ 423 ] = 32'h230FE040;
  assign memory[ 424 ] = 32'h2234446B;
  assign memory[ 425 ] = 32'hE03B701A;
  assign memory[ 426 ] = 32'h446B230F;
  assign memory[ 427 ] = 32'h701A2235;
  assign memory[ 428 ] = 32'h230FE036;
  assign memory[ 429 ] = 32'h2236446B;
  assign memory[ 430 ] = 32'hE031701A;
  assign memory[ 431 ] = 32'h446B230F;
  assign memory[ 432 ] = 32'h701A2237;
  assign memory[ 433 ] = 32'h230FE02C;
  assign memory[ 434 ] = 32'h2238446B;
  assign memory[ 435 ] = 32'hE027701A;
  assign memory[ 436 ] = 32'h446B230F;
  assign memory[ 437 ] = 32'h701A2239;
  assign memory[ 438 ] = 32'h230FE022;
  assign memory[ 439 ] = 32'h2241446B;
  assign memory[ 440 ] = 32'hE01D701A;
  assign memory[ 441 ] = 32'h446B230F;
  assign memory[ 442 ] = 32'h701A2242;
  assign memory[ 443 ] = 32'h230FE018;
  assign memory[ 444 ] = 32'h2243446B;
  assign memory[ 445 ] = 32'hE013701A;
  assign memory[ 446 ] = 32'h446B230F;
  assign memory[ 447 ] = 32'h701A2244;
  assign memory[ 448 ] = 32'h230FE00E;
  assign memory[ 449 ] = 32'h2245446B;
  assign memory[ 450 ] = 32'hE009701A;
  assign memory[ 451 ] = 32'h446B230F;
  assign memory[ 452 ] = 32'h701A2246;
  assign memory[ 453 ] = 32'h230FE004;
  assign memory[ 454 ] = 32'h2220446B;
  assign memory[ 455 ] = 32'h46C0701A;
  assign memory[ 456 ] = 32'h446B230F;
  assign memory[ 457 ] = 32'h0018781B;
  assign memory[ 458 ] = 32'h4770B004;
  assign memory[ 459 ] = 32'h000022D8;
  assign memory[ 460 ] = 32'hB08BB500;
  assign memory[ 461 ] = 32'h9B019001;
  assign memory[ 462 ] = 32'h0018494A;
  assign memory[ 463 ] = 32'hFB22F001;
  assign memory[ 464 ] = 32'h4949000B;
  assign memory[ 465 ] = 32'hF0010018;
  assign memory[ 466 ] = 32'h0003FA97;
  assign memory[ 467 ] = 32'h9B019309;
  assign memory[ 468 ] = 32'h00184945;
  assign memory[ 469 ] = 32'hFB16F001;
  assign memory[ 470 ] = 32'h4944000B;
  assign memory[ 471 ] = 32'hF0010018;
  assign memory[ 472 ] = 32'h0003FA8B;
  assign memory[ 473 ] = 32'h9B019308;
  assign memory[ 474 ] = 32'h00184940;
  assign memory[ 475 ] = 32'hFB0AF001;
  assign memory[ 476 ] = 32'h001A000B;
  assign memory[ 477 ] = 32'h009923FA;
  assign memory[ 478 ] = 32'hF0010010;
  assign memory[ 479 ] = 32'h0003FA7D;
  assign memory[ 480 ] = 32'h9A019307;
  assign memory[ 481 ] = 32'h009923FA;
  assign memory[ 482 ] = 32'hF0010010;
  assign memory[ 483 ] = 32'h000BFAFB;
  assign memory[ 484 ] = 32'h00182164;
  assign memory[ 485 ] = 32'hFA70F001;
  assign memory[ 486 ] = 32'h93060003;
  assign memory[ 487 ] = 32'h2B009B09;
  assign memory[ 488 ] = 32'h2310D10B;
  assign memory[ 489 ] = 32'h9B089309;
  assign memory[ 490 ] = 32'hD1062B00;
  assign memory[ 491 ] = 32'h93082310;
  assign memory[ 492 ] = 32'h2B009B07;
  assign memory[ 493 ] = 32'h2310D101;
  assign memory[ 494 ] = 32'hAB029307;
  assign memory[ 495 ] = 32'h701A2220;
  assign memory[ 496 ] = 32'h00189B09;
  assign memory[ 497 ] = 32'hFF4CF7FF;
  assign memory[ 498 ] = 32'h001A0003;
  assign memory[ 499 ] = 32'h705AAB02;
  assign memory[ 500 ] = 32'h00189B08;
  assign memory[ 501 ] = 32'hFF44F7FF;
  assign memory[ 502 ] = 32'h001A0003;
  assign memory[ 503 ] = 32'h709AAB02;
  assign memory[ 504 ] = 32'h00189B07;
  assign memory[ 505 ] = 32'hFF3CF7FF;
  assign memory[ 506 ] = 32'h001A0003;
  assign memory[ 507 ] = 32'h70DAAB02;
  assign memory[ 508 ] = 32'h00189B06;
  assign memory[ 509 ] = 32'hFF34F7FF;
  assign memory[ 510 ] = 32'h001A0003;
  assign memory[ 511 ] = 32'h711AAB02;
  assign memory[ 512 ] = 32'h2220AB02;
  assign memory[ 513 ] = 32'hAB02715A;
  assign memory[ 514 ] = 32'h719A226D;
  assign memory[ 515 ] = 32'h2262AB02;
  assign memory[ 516 ] = 32'hAB0271DA;
  assign memory[ 517 ] = 32'h061A79DB;
  assign memory[ 518 ] = 32'h799BAB02;
  assign memory[ 519 ] = 32'h18D2041B;
  assign memory[ 520 ] = 32'h795BAB02;
  assign memory[ 521 ] = 32'h18D3021B;
  assign memory[ 522 ] = 32'h7912AA02;
  assign memory[ 523 ] = 32'h9305189B;
  assign memory[ 524 ] = 32'h78DBAB02;
  assign memory[ 525 ] = 32'hAB02061A;
  assign memory[ 526 ] = 32'h041B789B;
  assign memory[ 527 ] = 32'hAB0218D2;
  assign memory[ 528 ] = 32'h021B785B;
  assign memory[ 529 ] = 32'hAA0218D3;
  assign memory[ 530 ] = 32'h189B7812;
  assign memory[ 531 ] = 32'h9B059304;
  assign memory[ 532 ] = 32'hF7FF0018;
  assign memory[ 533 ] = 32'h9B04FDC7;
  assign memory[ 534 ] = 32'hF7FF0018;
  assign memory[ 535 ] = 32'h46C0FDB7;
  assign memory[ 536 ] = 32'hBD00B00B;
  assign memory[ 537 ] = 32'h000F4240;
  assign memory[ 538 ] = 32'h000186A0;
  assign memory[ 539 ] = 32'h00002710;
  assign memory[ 540 ] = 32'hB08BB500;
  assign memory[ 541 ] = 32'h9B019001;
  assign memory[ 542 ] = 32'h00184948;
  assign memory[ 543 ] = 32'hFA82F001;
  assign memory[ 544 ] = 32'h001A000B;
  assign memory[ 545 ] = 32'h009923FA;
  assign memory[ 546 ] = 32'hF0010010;
  assign memory[ 547 ] = 32'h0003F9F5;
  assign memory[ 548 ] = 32'h9A019309;
  assign memory[ 549 ] = 32'h009923FA;
  assign memory[ 550 ] = 32'hF0010010;
  assign memory[ 551 ] = 32'h000BFA73;
  assign memory[ 552 ] = 32'h00182164;
  assign memory[ 553 ] = 32'hF9E8F001;
  assign memory[ 554 ] = 32'h93080003;
  assign memory[ 555 ] = 32'h21649B01;
  assign memory[ 556 ] = 32'hF0010018;
  assign memory[ 557 ] = 32'h000BFA67;
  assign memory[ 558 ] = 32'h0018210A;
  assign memory[ 559 ] = 32'hF9DCF001;
  assign memory[ 560 ] = 32'h93070003;
  assign memory[ 561 ] = 32'h210A9B01;
  assign memory[ 562 ] = 32'hF0010018;
  assign memory[ 563 ] = 32'h000BFA5B;
  assign memory[ 564 ] = 32'h9B099306;
  assign memory[ 565 ] = 32'hD10B2B00;
  assign memory[ 566 ] = 32'h93092310;
  assign memory[ 567 ] = 32'h2B009B08;
  assign memory[ 568 ] = 32'h2310D106;
  assign memory[ 569 ] = 32'h9B079308;
  assign memory[ 570 ] = 32'hD1012B00;
  assign memory[ 571 ] = 32'h93072310;
  assign memory[ 572 ] = 32'h2220AB02;
  assign memory[ 573 ] = 32'h9B09701A;
  assign memory[ 574 ] = 32'hF7FF0018;
  assign memory[ 575 ] = 32'h0003FEB1;
  assign memory[ 576 ] = 32'hAB02001A;
  assign memory[ 577 ] = 32'h9B08705A;
  assign memory[ 578 ] = 32'hF7FF0018;
  assign memory[ 579 ] = 32'h0003FEA9;
  assign memory[ 580 ] = 32'hAB02001A;
  assign memory[ 581 ] = 32'h9B07709A;
  assign memory[ 582 ] = 32'hF7FF0018;
  assign memory[ 583 ] = 32'h0003FEA1;
  assign memory[ 584 ] = 32'hAB02001A;
  assign memory[ 585 ] = 32'h9B0670DA;
  assign memory[ 586 ] = 32'hF7FF0018;
  assign memory[ 587 ] = 32'h0003FE99;
  assign memory[ 588 ] = 32'hAB02001A;
  assign memory[ 589 ] = 32'hAB02711A;
  assign memory[ 590 ] = 32'h715A2220;
  assign memory[ 591 ] = 32'h226DAB02;
  assign memory[ 592 ] = 32'hAB02719A;
  assign memory[ 593 ] = 32'h71DA2220;
  assign memory[ 594 ] = 32'h79DBAB02;
  assign memory[ 595 ] = 32'hAB02061A;
  assign memory[ 596 ] = 32'h041B799B;
  assign memory[ 597 ] = 32'hAB0218D2;
  assign memory[ 598 ] = 32'h021B795B;
  assign memory[ 599 ] = 32'hAA0218D3;
  assign memory[ 600 ] = 32'h189B7912;
  assign memory[ 601 ] = 32'hAB029305;
  assign memory[ 602 ] = 32'h061A78DB;
  assign memory[ 603 ] = 32'h789BAB02;
  assign memory[ 604 ] = 32'h18D2041B;
  assign memory[ 605 ] = 32'h785BAB02;
  assign memory[ 606 ] = 32'h18D3021B;
  assign memory[ 607 ] = 32'h7812AA02;
  assign memory[ 608 ] = 32'h9304189B;
  assign memory[ 609 ] = 32'h00189B05;
  assign memory[ 610 ] = 32'hFD2CF7FF;
  assign memory[ 611 ] = 32'h00189B04;
  assign memory[ 612 ] = 32'hFD1CF7FF;
  assign memory[ 613 ] = 32'hB00B46C0;
  assign memory[ 614 ] = 32'h46C0BD00;
  assign memory[ 615 ] = 32'h00002710;
  assign memory[ 616 ] = 32'hB08FB500;
  assign memory[ 617 ] = 32'h9A019001;
  assign memory[ 618 ] = 32'h011923E1;
  assign memory[ 619 ] = 32'hF0010010;
  assign memory[ 620 ] = 32'h0003F9ED;
  assign memory[ 621 ] = 32'h9A01930D;
  assign memory[ 622 ] = 32'h011923E1;
  assign memory[ 623 ] = 32'hF0010010;
  assign memory[ 624 ] = 32'h000BFACB;
  assign memory[ 625 ] = 32'h0018213C;
  assign memory[ 626 ] = 32'hF9E0F001;
  assign memory[ 627 ] = 32'h930C0003;
  assign memory[ 628 ] = 32'h213C9B01;
  assign memory[ 629 ] = 32'hF0010018;
  assign memory[ 630 ] = 32'h000BFABF;
  assign memory[ 631 ] = 32'h9B0D930B;
  assign memory[ 632 ] = 32'h0018210A;
  assign memory[ 633 ] = 32'hF9CEF001;
  assign memory[ 634 ] = 32'h930A000B;
  assign memory[ 635 ] = 32'h210A9B0C;
  assign memory[ 636 ] = 32'hF0010018;
  assign memory[ 637 ] = 32'h0003F941;
  assign memory[ 638 ] = 32'h9B0C9309;
  assign memory[ 639 ] = 32'h0018210A;
  assign memory[ 640 ] = 32'hF9C0F001;
  assign memory[ 641 ] = 32'h9308000B;
  assign memory[ 642 ] = 32'h210A9B0B;
  assign memory[ 643 ] = 32'hF0010018;
  assign memory[ 644 ] = 32'h0003F933;
  assign memory[ 645 ] = 32'h9B0B9307;
  assign memory[ 646 ] = 32'h0018210A;
  assign memory[ 647 ] = 32'hF9B2F001;
  assign memory[ 648 ] = 32'h9306000B;
  assign memory[ 649 ] = 32'h2220AB02;
  assign memory[ 650 ] = 32'h9B0A701A;
  assign memory[ 651 ] = 32'hF7FF0018;
  assign memory[ 652 ] = 32'h0003FE17;
  assign memory[ 653 ] = 32'hAB02001A;
  assign memory[ 654 ] = 32'hAB02705A;
  assign memory[ 655 ] = 32'h709A223A;
  assign memory[ 656 ] = 32'h00189B09;
  assign memory[ 657 ] = 32'hFE0CF7FF;
  assign memory[ 658 ] = 32'h001A0003;
  assign memory[ 659 ] = 32'h70DAAB02;
  assign memory[ 660 ] = 32'h00189B08;
  assign memory[ 661 ] = 32'hFE04F7FF;
  assign memory[ 662 ] = 32'h001A0003;
  assign memory[ 663 ] = 32'h711AAB02;
  assign memory[ 664 ] = 32'h223AAB02;
  assign memory[ 665 ] = 32'h9B07715A;
  assign memory[ 666 ] = 32'hF7FF0018;
  assign memory[ 667 ] = 32'h0003FDF9;
  assign memory[ 668 ] = 32'hAB02001A;
  assign memory[ 669 ] = 32'h9B06719A;
  assign memory[ 670 ] = 32'hF7FF0018;
  assign memory[ 671 ] = 32'h0003FDF1;
  assign memory[ 672 ] = 32'hAB02001A;
  assign memory[ 673 ] = 32'hAB0271DA;
  assign memory[ 674 ] = 32'h061A79DB;
  assign memory[ 675 ] = 32'h799BAB02;
  assign memory[ 676 ] = 32'h18D2041B;
  assign memory[ 677 ] = 32'h795BAB02;
  assign memory[ 678 ] = 32'h18D3021B;
  assign memory[ 679 ] = 32'h7912AA02;
  assign memory[ 680 ] = 32'h9305189B;
  assign memory[ 681 ] = 32'h78DBAB02;
  assign memory[ 682 ] = 32'hAB02061A;
  assign memory[ 683 ] = 32'h041B789B;
  assign memory[ 684 ] = 32'hAB0218D2;
  assign memory[ 685 ] = 32'h021B785B;
  assign memory[ 686 ] = 32'hAA0218D3;
  assign memory[ 687 ] = 32'h189B7812;
  assign memory[ 688 ] = 32'h9B059304;
  assign memory[ 689 ] = 32'hF7FF0018;
  assign memory[ 690 ] = 32'h9B04FC8D;
  assign memory[ 691 ] = 32'hF7FF0018;
  assign memory[ 692 ] = 32'h46C0FC7D;
  assign memory[ 693 ] = 32'hBD00B00F;
  assign memory[ 694 ] = 32'hB08DB500;
  assign memory[ 695 ] = 32'h9B019001;
  assign memory[ 696 ] = 32'h07DA0FDB;
  assign memory[ 697 ] = 32'h446B232B;
  assign memory[ 698 ] = 32'h418A1E51;
  assign memory[ 699 ] = 32'h9B01701A;
  assign memory[ 700 ] = 32'h232B930B;
  assign memory[ 701 ] = 32'h781B446B;
  assign memory[ 702 ] = 32'hD0022B00;
  assign memory[ 703 ] = 32'h425B9B0B;
  assign memory[ 704 ] = 32'h9B0B930B;
  assign memory[ 705 ] = 32'h210A139B;
  assign memory[ 706 ] = 32'hF0010018;
  assign memory[ 707 ] = 32'h000BFA25;
  assign memory[ 708 ] = 32'h9A0B9309;
  assign memory[ 709 ] = 32'h009B0013;
  assign memory[ 710 ] = 32'h005B189B;
  assign memory[ 711 ] = 32'h210A139B;
  assign memory[ 712 ] = 32'hF0010018;
  assign memory[ 713 ] = 32'h000BFA19;
  assign memory[ 714 ] = 32'h9B0B9308;
  assign memory[ 715 ] = 32'h43532264;
  assign memory[ 716 ] = 32'h210A139B;
  assign memory[ 717 ] = 32'hF0010018;
  assign memory[ 718 ] = 32'h000BFA0F;
  assign memory[ 719 ] = 32'h232B9307;
  assign memory[ 720 ] = 32'h781B446B;
  assign memory[ 721 ] = 32'hD0032B00;
  assign memory[ 722 ] = 32'h222DAB03;
  assign memory[ 723 ] = 32'hE002701A;
  assign memory[ 724 ] = 32'h2220AB03;
  assign memory[ 725 ] = 32'h9B09701A;
  assign memory[ 726 ] = 32'hF7FF0018;
  assign memory[ 727 ] = 32'h0003FD81;
  assign memory[ 728 ] = 32'hAB03001A;
  assign memory[ 729 ] = 32'hAB03705A;
  assign memory[ 730 ] = 32'h709A222E;
  assign memory[ 731 ] = 32'h00189B08;
  assign memory[ 732 ] = 32'hFD76F7FF;
  assign memory[ 733 ] = 32'h001A0003;
  assign memory[ 734 ] = 32'h70DAAB03;
  assign memory[ 735 ] = 32'h00189B07;
  assign memory[ 736 ] = 32'hFD6EF7FF;
  assign memory[ 737 ] = 32'h001A0003;
  assign memory[ 738 ] = 32'h711AAB03;
  assign memory[ 739 ] = 32'h226DAB03;
  assign memory[ 740 ] = 32'hAB03715A;
  assign memory[ 741 ] = 32'h719A222F;
  assign memory[ 742 ] = 32'h2273AB03;
  assign memory[ 743 ] = 32'hAB0371DA;
  assign memory[ 744 ] = 32'h061A79DB;
  assign memory[ 745 ] = 32'h799BAB03;
  assign memory[ 746 ] = 32'h18D2041B;
  assign memory[ 747 ] = 32'h795BAB03;
  assign memory[ 748 ] = 32'h18D3021B;
  assign memory[ 749 ] = 32'h7912AA03;
  assign memory[ 750 ] = 32'h9306189B;
  assign memory[ 751 ] = 32'h78DBAB03;
  assign memory[ 752 ] = 32'hAB03061A;
  assign memory[ 753 ] = 32'h041B789B;
  assign memory[ 754 ] = 32'hAB0318D2;
  assign memory[ 755 ] = 32'h021B785B;
  assign memory[ 756 ] = 32'hAA0318D3;
  assign memory[ 757 ] = 32'h189B7812;
  assign memory[ 758 ] = 32'h9B069305;
  assign memory[ 759 ] = 32'hF7FF0018;
  assign memory[ 760 ] = 32'h9B05FC01;
  assign memory[ 761 ] = 32'hF7FF0018;
  assign memory[ 762 ] = 32'h46C0FBF1;
  assign memory[ 763 ] = 32'hBD00B00D;
  assign memory[ 764 ] = 32'hB087B500;
  assign memory[ 765 ] = 32'h9B019001;
  assign memory[ 766 ] = 32'h781B3305;
  assign memory[ 767 ] = 32'hF7FF0018;
  assign memory[ 768 ] = 32'h0003FD2F;
  assign memory[ 769 ] = 32'hAB02001A;
  assign memory[ 770 ] = 32'h9B01701A;
  assign memory[ 771 ] = 32'h781B3304;
  assign memory[ 772 ] = 32'hF7FF0018;
  assign memory[ 773 ] = 32'h0003FD25;
  assign memory[ 774 ] = 32'hAB02001A;
  assign memory[ 775 ] = 32'h9B01705A;
  assign memory[ 776 ] = 32'h781B3303;
  assign memory[ 777 ] = 32'hF7FF0018;
  assign memory[ 778 ] = 32'h0003FD1B;
  assign memory[ 779 ] = 32'hAB02001A;
  assign memory[ 780 ] = 32'h9B01709A;
  assign memory[ 781 ] = 32'h781B3302;
  assign memory[ 782 ] = 32'hF7FF0018;
  assign memory[ 783 ] = 32'h0003FD11;
  assign memory[ 784 ] = 32'hAB02001A;
  assign memory[ 785 ] = 32'h9B0170DA;
  assign memory[ 786 ] = 32'h781B3301;
  assign memory[ 787 ] = 32'hF7FF0018;
  assign memory[ 788 ] = 32'h0003FD07;
  assign memory[ 789 ] = 32'hAB02001A;
  assign memory[ 790 ] = 32'h9B01711A;
  assign memory[ 791 ] = 32'h0018781B;
  assign memory[ 792 ] = 32'hFCFEF7FF;
  assign memory[ 793 ] = 32'h001A0003;
  assign memory[ 794 ] = 32'h715AAB02;
  assign memory[ 795 ] = 32'h2250AB02;
  assign memory[ 796 ] = 32'hAB02719A;
  assign memory[ 797 ] = 32'h71DA2261;
  assign memory[ 798 ] = 32'h79DBAB02;
  assign memory[ 799 ] = 32'hAB02061A;
  assign memory[ 800 ] = 32'h041B799B;
  assign memory[ 801 ] = 32'hAB0218D2;
  assign memory[ 802 ] = 32'h021B795B;
  assign memory[ 803 ] = 32'hAA0218D3;
  assign memory[ 804 ] = 32'h189B7912;
  assign memory[ 805 ] = 32'hAB029305;
  assign memory[ 806 ] = 32'h061A78DB;
  assign memory[ 807 ] = 32'h789BAB02;
  assign memory[ 808 ] = 32'h18D2041B;
  assign memory[ 809 ] = 32'h785BAB02;
  assign memory[ 810 ] = 32'h18D3021B;
  assign memory[ 811 ] = 32'h7812AA02;
  assign memory[ 812 ] = 32'h9304189B;
  assign memory[ 813 ] = 32'h00189B05;
  assign memory[ 814 ] = 32'hFB94F7FF;
  assign memory[ 815 ] = 32'h00189B04;
  assign memory[ 816 ] = 32'hFB84F7FF;
  assign memory[ 817 ] = 32'hB00746C0;
  assign memory[ 818 ] = 32'h46C0BD00;
  assign memory[ 819 ] = 32'hB087B500;
  assign memory[ 820 ] = 32'hAB029001;
  assign memory[ 821 ] = 32'h701A2220;
  assign memory[ 822 ] = 32'h33039B01;
  assign memory[ 823 ] = 32'h0018781B;
  assign memory[ 824 ] = 32'hFCBEF7FF;
  assign memory[ 825 ] = 32'h001A0003;
  assign memory[ 826 ] = 32'h705AAB02;
  assign memory[ 827 ] = 32'h33029B01;
  assign memory[ 828 ] = 32'h0018781B;
  assign memory[ 829 ] = 32'hFCB4F7FF;
  assign memory[ 830 ] = 32'h001A0003;
  assign memory[ 831 ] = 32'h709AAB02;
  assign memory[ 832 ] = 32'h33019B01;
  assign memory[ 833 ] = 32'h0018781B;
  assign memory[ 834 ] = 32'hFCAAF7FF;
  assign memory[ 835 ] = 32'h001A0003;
  assign memory[ 836 ] = 32'h70DAAB02;
  assign memory[ 837 ] = 32'h781B9B01;
  assign memory[ 838 ] = 32'hF7FF0018;
  assign memory[ 839 ] = 32'h0003FCA1;
  assign memory[ 840 ] = 32'hAB02001A;
  assign memory[ 841 ] = 32'hAB02711A;
  assign memory[ 842 ] = 32'h715A2220;
  assign memory[ 843 ] = 32'h226DAB02;
  assign memory[ 844 ] = 32'hAB02719A;
  assign memory[ 845 ] = 32'h71DA2220;
  assign memory[ 846 ] = 32'h79DBAB02;
  assign memory[ 847 ] = 32'hAB02061A;
  assign memory[ 848 ] = 32'h041B799B;
  assign memory[ 849 ] = 32'hAB0218D2;
  assign memory[ 850 ] = 32'h021B795B;
  assign memory[ 851 ] = 32'hAA0218D3;
  assign memory[ 852 ] = 32'h189B7912;
  assign memory[ 853 ] = 32'hAB029305;
  assign memory[ 854 ] = 32'h061A78DB;
  assign memory[ 855 ] = 32'h789BAB02;
  assign memory[ 856 ] = 32'h18D2041B;
  assign memory[ 857 ] = 32'h785BAB02;
  assign memory[ 858 ] = 32'h18D3021B;
  assign memory[ 859 ] = 32'h7812AA02;
  assign memory[ 860 ] = 32'h9304189B;
  assign memory[ 861 ] = 32'h00189B05;
  assign memory[ 862 ] = 32'hFB34F7FF;
  assign memory[ 863 ] = 32'h00189B04;
  assign memory[ 864 ] = 32'hFB24F7FF;
  assign memory[ 865 ] = 32'hB00746C0;
  assign memory[ 866 ] = 32'h46C0BD00;
  assign memory[ 867 ] = 32'h231BB510;
  assign memory[ 868 ] = 32'h211D221C;
  assign memory[ 869 ] = 32'hF7FF2000;
  assign memory[ 870 ] = 32'h2333FA77;
  assign memory[ 871 ] = 32'h21022202;
  assign memory[ 872 ] = 32'hF7FF2000;
  assign memory[ 873 ] = 32'h2103FAC5;
  assign memory[ 874 ] = 32'hF7FF2000;
  assign memory[ 875 ] = 32'h46C0FAF5;
  assign memory[ 876 ] = 32'hFA48F7FF;
  assign memory[ 877 ] = 32'hD1FB1E03;
  assign memory[ 878 ] = 32'hBD1046C0;
  assign memory[ 879 ] = 32'hB089B500;
  assign memory[ 880 ] = 32'h00119100;
  assign memory[ 881 ] = 32'h3307466B;
  assign memory[ 882 ] = 32'h701A1C02;
  assign memory[ 883 ] = 32'h3306466B;
  assign memory[ 884 ] = 32'h701A1C0A;
  assign memory[ 885 ] = 32'h3307466B;
  assign memory[ 886 ] = 32'h2200781B;
  assign memory[ 887 ] = 32'h20002100;
  assign memory[ 888 ] = 32'hFA52F7FF;
  assign memory[ 889 ] = 32'hF7FF46C0;
  assign memory[ 890 ] = 32'h1E03FA2D;
  assign memory[ 891 ] = 32'h466BD1FB;
  assign memory[ 892 ] = 32'h781B3306;
  assign memory[ 893 ] = 32'h20010019;
  assign memory[ 894 ] = 32'hFACEF7FF;
  assign memory[ 895 ] = 32'hF7FF46C0;
  assign memory[ 896 ] = 32'h0003FA13;
  assign memory[ 897 ] = 32'h2301001A;
  assign memory[ 898 ] = 32'hB2DB4053;
  assign memory[ 899 ] = 32'hD1F62B00;
  assign memory[ 900 ] = 32'h3306466B;
  assign memory[ 901 ] = 32'h2B03781B;
  assign memory[ 902 ] = 32'hF7FFD822;
  assign memory[ 903 ] = 32'h0003FA71;
  assign memory[ 904 ] = 32'h23FF9306;
  assign memory[ 905 ] = 32'h23009305;
  assign memory[ 906 ] = 32'hE0129307;
  assign memory[ 907 ] = 32'h9B079A00;
  assign memory[ 908 ] = 32'h9A0718D3;
  assign memory[ 909 ] = 32'h990500D2;
  assign memory[ 910 ] = 32'h000A4091;
  assign memory[ 911 ] = 32'h40119906;
  assign memory[ 912 ] = 32'h00D29A07;
  assign memory[ 913 ] = 32'h000A40D1;
  assign memory[ 914 ] = 32'h701AB2D2;
  assign memory[ 915 ] = 32'h33019B07;
  assign memory[ 916 ] = 32'h466B9307;
  assign memory[ 917 ] = 32'h781A3306;
  assign memory[ 918 ] = 32'h429A9B07;
  assign memory[ 919 ] = 32'hE03FD8E6;
  assign memory[ 920 ] = 32'hFA4EF7FF;
  assign memory[ 921 ] = 32'h93060003;
  assign memory[ 922 ] = 32'hFA52F7FF;
  assign memory[ 923 ] = 32'h93040003;
  assign memory[ 924 ] = 32'h930323FF;
  assign memory[ 925 ] = 32'h93072300;
  assign memory[ 926 ] = 32'h9B07E02C;
  assign memory[ 927 ] = 32'hD8102B03;
  assign memory[ 928 ] = 32'h9B079A00;
  assign memory[ 929 ] = 32'h9A0718D3;
  assign memory[ 930 ] = 32'h990300D2;
  assign memory[ 931 ] = 32'h000A4091;
  assign memory[ 932 ] = 32'h40119906;
  assign memory[ 933 ] = 32'h00D29A07;
  assign memory[ 934 ] = 32'h000A40D1;
  assign memory[ 935 ] = 32'h701AB2D2;
  assign memory[ 936 ] = 32'h9A00E015;
  assign memory[ 937 ] = 32'h18D39B07;
  assign memory[ 938 ] = 32'h490F9A07;
  assign memory[ 939 ] = 32'h4462468C;
  assign memory[ 940 ] = 32'h990300D2;
  assign memory[ 941 ] = 32'h000A4091;
  assign memory[ 942 ] = 32'h40119904;
  assign memory[ 943 ] = 32'h480A9A07;
  assign memory[ 944 ] = 32'h44624684;
  assign memory[ 945 ] = 32'h40D100D2;
  assign memory[ 946 ] = 32'hB2D2000A;
  assign memory[ 947 ] = 32'h9B07701A;
  assign memory[ 948 ] = 32'h93073301;
  assign memory[ 949 ] = 32'h3306466B;
  assign memory[ 950 ] = 32'h9B07781A;
  assign memory[ 951 ] = 32'hD8CC429A;
  assign memory[ 952 ] = 32'hB00946C0;
  assign memory[ 953 ] = 32'h46C0BD00;
  assign memory[ 954 ] = 32'h1FFFFFFC;
  assign memory[ 955 ] = 32'hB085B500;
  assign memory[ 956 ] = 32'hAB029001;
  assign memory[ 957 ] = 32'h00192205;
  assign memory[ 958 ] = 32'hF7FF2031;
  assign memory[ 959 ] = 32'hAB02FF5F;
  assign memory[ 960 ] = 32'h021B785B;
  assign memory[ 961 ] = 32'hAB02B21A;
  assign memory[ 962 ] = 32'hB21B781B;
  assign memory[ 963 ] = 32'hB21B4313;
  assign memory[ 964 ] = 32'h9B01B29A;
  assign memory[ 965 ] = 32'hAB02801A;
  assign memory[ 966 ] = 32'h021B78DB;
  assign memory[ 967 ] = 32'hAB02B21A;
  assign memory[ 968 ] = 32'hB21B789B;
  assign memory[ 969 ] = 32'hB21B4313;
  assign memory[ 970 ] = 32'h9B01B29A;
  assign memory[ 971 ] = 32'hAB02805A;
  assign memory[ 972 ] = 32'hB25A791B;
  assign memory[ 973 ] = 32'h711A9B01;
  assign memory[ 974 ] = 32'h2206AB02;
  assign memory[ 975 ] = 32'h20360019;
  assign memory[ 976 ] = 32'hFF3CF7FF;
  assign memory[ 977 ] = 32'h785BAB02;
  assign memory[ 978 ] = 32'hB21A021B;
  assign memory[ 979 ] = 32'h781BAB02;
  assign memory[ 980 ] = 32'h4313B21B;
  assign memory[ 981 ] = 32'h9B01B21A;
  assign memory[ 982 ] = 32'hAB0280DA;
  assign memory[ 983 ] = 32'h021B78DB;
  assign memory[ 984 ] = 32'hAB02B21A;
  assign memory[ 985 ] = 32'hB21B789B;
  assign memory[ 986 ] = 32'hB21A4313;
  assign memory[ 987 ] = 32'h811A9B01;
  assign memory[ 988 ] = 32'h791BAB02;
  assign memory[ 989 ] = 32'h9B01B25A;
  assign memory[ 990 ] = 32'hAB02729A;
  assign memory[ 991 ] = 32'hB25A795B;
  assign memory[ 992 ] = 32'h72DA9B01;
  assign memory[ 993 ] = 32'h2206AB02;
  assign memory[ 994 ] = 32'h203C0019;
  assign memory[ 995 ] = 32'hFF16F7FF;
  assign memory[ 996 ] = 32'h785BAB02;
  assign memory[ 997 ] = 32'hB21A021B;
  assign memory[ 998 ] = 32'h781BAB02;
  assign memory[ 999 ] = 32'h4313B21B;
  assign memory[ 1000 ] = 32'hB29AB21B;
  assign memory[ 1001 ] = 32'h819A9B01;
  assign memory[ 1002 ] = 32'h78DBAB02;
  assign memory[ 1003 ] = 32'hB21A021B;
  assign memory[ 1004 ] = 32'h789BAB02;
  assign memory[ 1005 ] = 32'h4313B21B;
  assign memory[ 1006 ] = 32'hB29AB21B;
  assign memory[ 1007 ] = 32'h81DA9B01;
  assign memory[ 1008 ] = 32'h791BAB02;
  assign memory[ 1009 ] = 32'h9B01B25A;
  assign memory[ 1010 ] = 32'hAB02741A;
  assign memory[ 1011 ] = 32'hB25A795B;
  assign memory[ 1012 ] = 32'h745A9B01;
  assign memory[ 1013 ] = 32'h2204AB02;
  assign memory[ 1014 ] = 32'h20420019;
  assign memory[ 1015 ] = 32'hFEEEF7FF;
  assign memory[ 1016 ] = 32'h785BAB02;
  assign memory[ 1017 ] = 32'hB21A021B;
  assign memory[ 1018 ] = 32'h781BAB02;
  assign memory[ 1019 ] = 32'h4313B21B;
  assign memory[ 1020 ] = 32'h9B01B21A;
  assign memory[ 1021 ] = 32'hAB02825A;
  assign memory[ 1022 ] = 32'hB25A789B;
  assign memory[ 1023 ] = 32'h751A9B01;
  assign memory[ 1024 ] = 32'h78DBAB02;
  assign memory[ 1025 ] = 32'h9B01B25A;
  assign memory[ 1026 ] = 32'h46C0755A;
  assign memory[ 1027 ] = 32'hBD00B005;
  assign memory[ 1028 ] = 32'hB099B5F0;
  assign memory[ 1029 ] = 32'h91089009;
  assign memory[ 1030 ] = 32'h92009A09;
  assign memory[ 1031 ] = 32'h92012200;
  assign memory[ 1032 ] = 32'h88129A08;
  assign memory[ 1033 ] = 32'h22009202;
  assign memory[ 1034 ] = 32'h98029203;
  assign memory[ 1035 ] = 32'h00029903;
  assign memory[ 1036 ] = 32'h000F0E12;
  assign memory[ 1037 ] = 32'h4314023C;
  assign memory[ 1038 ] = 32'h02130002;
  assign memory[ 1039 ] = 32'h9A019900;
  assign memory[ 1040 ] = 32'h41A21AC9;
  assign memory[ 1041 ] = 32'h0014000B;
  assign memory[ 1042 ] = 32'h94179316;
  assign memory[ 1043 ] = 32'h885B9B08;
  assign memory[ 1044 ] = 32'h23009304;
  assign memory[ 1045 ] = 32'h9A169305;
  assign memory[ 1046 ] = 32'h98049B17;
  assign memory[ 1047 ] = 32'hF0009905;
  assign memory[ 1048 ] = 32'h0003FFA5;
  assign memory[ 1049 ] = 32'h9314000C;
  assign memory[ 1050 ] = 32'h9A169415;
  assign memory[ 1051 ] = 32'h98169B17;
  assign memory[ 1052 ] = 32'hF0009917;
  assign memory[ 1053 ] = 32'h0003FF9B;
  assign memory[ 1054 ] = 32'h9312000C;
  assign memory[ 1055 ] = 32'h9B089413;
  assign memory[ 1056 ] = 32'hB25B791B;
  assign memory[ 1057 ] = 32'h17DB9306;
  assign memory[ 1058 ] = 32'h9B129307;
  assign memory[ 1059 ] = 32'h001A9C13;
  assign memory[ 1060 ] = 32'h98060023;
  assign memory[ 1061 ] = 32'hF0009907;
  assign memory[ 1062 ] = 32'h0003FF89;
  assign memory[ 1063 ] = 32'h9310000C;
  assign memory[ 1064 ] = 32'h9B149411;
  assign memory[ 1065 ] = 32'h0B9A9C15;
  assign memory[ 1066 ] = 32'h431604A6;
  assign memory[ 1067 ] = 32'h9B10049D;
  assign memory[ 1068 ] = 32'h195B9C11;
  assign memory[ 1069 ] = 32'h930E4174;
  assign memory[ 1070 ] = 32'h9B0F940F;
  assign memory[ 1071 ] = 32'h930C001B;
  assign memory[ 1072 ] = 32'h17DB9B0F;
  assign memory[ 1073 ] = 32'h9A08930D;
  assign memory[ 1074 ] = 32'h9C0D9B0C;
  assign memory[ 1075 ] = 32'h61D46193;
  assign memory[ 1076 ] = 32'h041B9B0D;
  assign memory[ 1077 ] = 32'h0C129A0C;
  assign memory[ 1078 ] = 32'h930A4313;
  assign memory[ 1079 ] = 32'h141B9B0D;
  assign memory[ 1080 ] = 32'h9B0A930B;
  assign memory[ 1081 ] = 32'h00189C0B;
  assign memory[ 1082 ] = 32'hB0190021;
  assign memory[ 1083 ] = 32'h46C0BDF0;
  assign memory[ 1084 ] = 32'hB0C0B570;
  assign memory[ 1085 ] = 32'h912C902D;
  assign memory[ 1086 ] = 32'h69989B2C;
  assign memory[ 1087 ] = 32'h9B2C69D9;
  assign memory[ 1088 ] = 32'h699B69DC;
  assign memory[ 1089 ] = 32'h0023001A;
  assign memory[ 1090 ] = 32'hFF50F000;
  assign memory[ 1091 ] = 32'h000C0003;
  assign memory[ 1092 ] = 32'h943F933E;
  assign memory[ 1093 ] = 32'h069A9B3F;
  assign memory[ 1094 ] = 32'h099B9B3E;
  assign memory[ 1095 ] = 32'h933C4313;
  assign memory[ 1096 ] = 32'h119B9B3F;
  assign memory[ 1097 ] = 32'h9B2C933D;
  assign memory[ 1098 ] = 32'h69D96998;
  assign memory[ 1099 ] = 32'h9B3D9A3C;
  assign memory[ 1100 ] = 32'hFF3CF000;
  assign memory[ 1101 ] = 32'h000C0003;
  assign memory[ 1102 ] = 32'h0A1A0621;
  assign memory[ 1103 ] = 32'h923A430A;
  assign memory[ 1104 ] = 32'h933B1223;
  assign memory[ 1105 ] = 32'h7C5B9B2C;
  assign memory[ 1106 ] = 32'h9306B25B;
  assign memory[ 1107 ] = 32'h930717DB;
  assign memory[ 1108 ] = 32'h9B3B9A3A;
  assign memory[ 1109 ] = 32'h99079806;
  assign memory[ 1110 ] = 32'hFF28F000;
  assign memory[ 1111 ] = 32'h000C0003;
  assign memory[ 1112 ] = 32'h095A06E1;
  assign memory[ 1113 ] = 32'h9238430A;
  assign memory[ 1114 ] = 32'h93391163;
  assign memory[ 1115 ] = 32'h7C1B9B2C;
  assign memory[ 1116 ] = 32'h9308B25B;
  assign memory[ 1117 ] = 32'h930917DB;
  assign memory[ 1118 ] = 32'h9B3F9A3E;
  assign memory[ 1119 ] = 32'h99099808;
  assign memory[ 1120 ] = 32'hFF14F000;
  assign memory[ 1121 ] = 32'h000C0003;
  assign memory[ 1122 ] = 32'h01220F19;
  assign memory[ 1123 ] = 32'h9237430A;
  assign memory[ 1124 ] = 32'h9336011B;
  assign memory[ 1125 ] = 32'h89DB9B2C;
  assign memory[ 1126 ] = 32'h2300930A;
  assign memory[ 1127 ] = 32'h9B2C930B;
  assign memory[ 1128 ] = 32'h699B69DC;
  assign memory[ 1129 ] = 32'h0023001A;
  assign memory[ 1130 ] = 32'h990B980A;
  assign memory[ 1131 ] = 32'hFEFEF000;
  assign memory[ 1132 ] = 32'h000C0003;
  assign memory[ 1133 ] = 32'h05A20A99;
  assign memory[ 1134 ] = 32'h9235430A;
  assign memory[ 1135 ] = 32'h9334059B;
  assign memory[ 1136 ] = 32'h899B9B2C;
  assign memory[ 1137 ] = 32'h2300930C;
  assign memory[ 1138 ] = 32'h9B0C930D;
  assign memory[ 1139 ] = 32'h930F03DB;
  assign memory[ 1140 ] = 32'h930E2300;
  assign memory[ 1141 ] = 32'h9C399B38;
  assign memory[ 1142 ] = 32'h9A0F990E;
  assign memory[ 1143 ] = 32'h416218C9;
  assign memory[ 1144 ] = 32'h9C379B36;
  assign memory[ 1145 ] = 32'h416218C9;
  assign memory[ 1146 ] = 32'h9C359B34;
  assign memory[ 1147 ] = 32'h4154185B;
  assign memory[ 1148 ] = 32'h94339332;
  assign memory[ 1149 ] = 32'h7ADB9B2C;
  assign memory[ 1150 ] = 32'h9310B25B;
  assign memory[ 1151 ] = 32'h931117DB;
  assign memory[ 1152 ] = 32'h9B3B9A3A;
  assign memory[ 1153 ] = 32'h99119810;
  assign memory[ 1154 ] = 32'hFED0F000;
  assign memory[ 1155 ] = 32'h000C0003;
  assign memory[ 1156 ] = 32'h095A06E1;
  assign memory[ 1157 ] = 32'h923C430A;
  assign memory[ 1158 ] = 32'h933D1163;
  assign memory[ 1159 ] = 32'h7A9B9B2C;
  assign memory[ 1160 ] = 32'h9312B25B;
  assign memory[ 1161 ] = 32'h931317DB;
  assign memory[ 1162 ] = 32'h9B3F9A3E;
  assign memory[ 1163 ] = 32'h99139812;
  assign memory[ 1164 ] = 32'hFEBCF000;
  assign memory[ 1165 ] = 32'h000C0003;
  assign memory[ 1166 ] = 32'h00A20F99;
  assign memory[ 1167 ] = 32'h9239430A;
  assign memory[ 1168 ] = 32'h9338009B;
  assign memory[ 1169 ] = 32'h22089B2C;
  assign memory[ 1170 ] = 32'h93145E9B;
  assign memory[ 1171 ] = 32'h931517DB;
  assign memory[ 1172 ] = 32'h24014B8C;
  assign memory[ 1173 ] = 32'h98144264;
  assign memory[ 1174 ] = 32'h18C09915;
  assign memory[ 1175 ] = 32'h9B2C4161;
  assign memory[ 1176 ] = 32'h699B69DC;
  assign memory[ 1177 ] = 32'h0023001A;
  assign memory[ 1178 ] = 32'hFEA0F000;
  assign memory[ 1179 ] = 32'h000C0003;
  assign memory[ 1180 ] = 32'h05620AD9;
  assign memory[ 1181 ] = 32'h9237430A;
  assign memory[ 1182 ] = 32'h9336055B;
  assign memory[ 1183 ] = 32'h22069B2C;
  assign memory[ 1184 ] = 32'h93165E9B;
  assign memory[ 1185 ] = 32'h931717DB;
  assign memory[ 1186 ] = 32'h24014B7E;
  assign memory[ 1187 ] = 32'h99164264;
  assign memory[ 1188 ] = 32'h18C99A17;
  assign memory[ 1189 ] = 32'h000B4162;
  assign memory[ 1190 ] = 32'h039B0014;
  assign memory[ 1191 ] = 32'h23009319;
  assign memory[ 1192 ] = 32'h9B3C9318;
  assign memory[ 1193 ] = 32'h99189C3D;
  assign memory[ 1194 ] = 32'h18C99A19;
  assign memory[ 1195 ] = 32'h9B384162;
  assign memory[ 1196 ] = 32'h18C99C39;
  assign memory[ 1197 ] = 32'h9B364162;
  assign memory[ 1198 ] = 32'h185B9C37;
  assign memory[ 1199 ] = 32'h93304154;
  assign memory[ 1200 ] = 32'h9B319431;
  assign memory[ 1201 ] = 32'h9B30021A;
  assign memory[ 1202 ] = 32'h93000E1B;
  assign memory[ 1203 ] = 32'h43139B00;
  assign memory[ 1204 ] = 32'h9B319300;
  assign memory[ 1205 ] = 32'h9301161B;
  assign memory[ 1206 ] = 32'h931A9B2D;
  assign memory[ 1207 ] = 32'h931B2300;
  assign memory[ 1208 ] = 32'h9B1B9A1A;
  assign memory[ 1209 ] = 32'h99019800;
  assign memory[ 1210 ] = 32'hFE60F000;
  assign memory[ 1211 ] = 32'h000C0003;
  assign memory[ 1212 ] = 32'h943F933E;
  assign memory[ 1213 ] = 32'h7D1B9B2C;
  assign memory[ 1214 ] = 32'h931CB25B;
  assign memory[ 1215 ] = 32'h931D17DB;
  assign memory[ 1216 ] = 32'h69DC9B2C;
  assign memory[ 1217 ] = 32'h001A699B;
  assign memory[ 1218 ] = 32'h981C0023;
  assign memory[ 1219 ] = 32'hF000991D;
  assign memory[ 1220 ] = 32'h0003FE4D;
  assign memory[ 1221 ] = 32'h933C000C;
  assign memory[ 1222 ] = 32'h9B2C943D;
  assign memory[ 1223 ] = 32'h5E9B2212;
  assign memory[ 1224 ] = 32'h17DB931E;
  assign memory[ 1225 ] = 32'h991E931F;
  assign memory[ 1226 ] = 32'h000B9A1F;
  assign memory[ 1227 ] = 32'h00100C1B;
  assign memory[ 1228 ] = 32'h431E0406;
  assign memory[ 1229 ] = 32'h041D000B;
  assign memory[ 1230 ] = 32'h9C3D9B3C;
  assign memory[ 1231 ] = 32'h4174195B;
  assign memory[ 1232 ] = 32'h943B933A;
  assign memory[ 1233 ] = 32'h93209B2D;
  assign memory[ 1234 ] = 32'h93212300;
  assign memory[ 1235 ] = 32'h9B3B9A3A;
  assign memory[ 1236 ] = 32'h99219820;
  assign memory[ 1237 ] = 32'hFE2AF000;
  assign memory[ 1238 ] = 32'h000C0003;
  assign memory[ 1239 ] = 32'h0B5A04E1;
  assign memory[ 1240 ] = 32'h9238430A;
  assign memory[ 1241 ] = 32'h93391363;
  assign memory[ 1242 ] = 32'h99399838;
  assign memory[ 1243 ] = 32'h2300220A;
  assign memory[ 1244 ] = 32'hFDF8F000;
  assign memory[ 1245 ] = 32'h000C0003;
  assign memory[ 1246 ] = 32'h00210018;
  assign memory[ 1247 ] = 32'h93229B2D;
  assign memory[ 1248 ] = 32'h93232300;
  assign memory[ 1249 ] = 32'h9B239A22;
  assign memory[ 1250 ] = 32'hFE10F000;
  assign memory[ 1251 ] = 32'h000C0003;
  assign memory[ 1252 ] = 32'h0A5A05E1;
  assign memory[ 1253 ] = 32'h9236430A;
  assign memory[ 1254 ] = 32'h93371263;
  assign memory[ 1255 ] = 32'h9A379936;
  assign memory[ 1256 ] = 32'h0014000B;
  assign memory[ 1257 ] = 32'h00A50F98;
  assign memory[ 1258 ] = 32'h9D059505;
  assign memory[ 1259 ] = 32'h95054305;
  assign memory[ 1260 ] = 32'h9304009B;
  assign memory[ 1261 ] = 32'h9C059B04;
  assign memory[ 1262 ] = 32'h4154185B;
  assign memory[ 1263 ] = 32'h416418DB;
  assign memory[ 1264 ] = 32'h94379336;
  assign memory[ 1265 ] = 32'h93249B2D;
  assign memory[ 1266 ] = 32'h93252300;
  assign memory[ 1267 ] = 32'h93269B2D;
  assign memory[ 1268 ] = 32'h93272300;
  assign memory[ 1269 ] = 32'h9B279A26;
  assign memory[ 1270 ] = 32'h99259824;
  assign memory[ 1271 ] = 32'hFDE6F000;
  assign memory[ 1272 ] = 32'h000C0003;
  assign memory[ 1273 ] = 32'h94359334;
  assign memory[ 1274 ] = 32'h7D5B9B2C;
  assign memory[ 1275 ] = 32'h9328B25B;
  assign memory[ 1276 ] = 32'h932917DB;
  assign memory[ 1277 ] = 32'h9B359A34;
  assign memory[ 1278 ] = 32'h99299828;
  assign memory[ 1279 ] = 32'hFDD6F000;
  assign memory[ 1280 ] = 32'h000C0003;
  assign memory[ 1281 ] = 32'h0C190422;
  assign memory[ 1282 ] = 32'h923C430A;
  assign memory[ 1283 ] = 32'h933D1423;
  assign memory[ 1284 ] = 32'h932A9B2D;
  assign memory[ 1285 ] = 32'h932B2300;
  assign memory[ 1286 ] = 32'h9B3D9A3C;
  assign memory[ 1287 ] = 32'h992B982A;
  assign memory[ 1288 ] = 32'hFDC4F000;
  assign memory[ 1289 ] = 32'h000C0003;
  assign memory[ 1290 ] = 32'h09D90662;
  assign memory[ 1291 ] = 32'h923A430A;
  assign memory[ 1292 ] = 32'h933B11E3;
  assign memory[ 1293 ] = 32'h079B9B33;
  assign memory[ 1294 ] = 32'h08929A32;
  assign memory[ 1295 ] = 32'h9A029202;
  assign memory[ 1296 ] = 32'h9202431A;
  assign memory[ 1297 ] = 32'h109B9B33;
  assign memory[ 1298 ] = 32'h9B3E9303;
  assign memory[ 1299 ] = 32'h99029C3F;
  assign memory[ 1300 ] = 32'h18C99A03;
  assign memory[ 1301 ] = 32'h9B364162;
  assign memory[ 1302 ] = 32'h18C99C37;
  assign memory[ 1303 ] = 32'h9B3A4162;
  assign memory[ 1304 ] = 32'h185B9C3B;
  assign memory[ 1305 ] = 32'h93384154;
  assign memory[ 1306 ] = 32'h9B389439;
  assign memory[ 1307 ] = 32'h0AA39C39;
  assign memory[ 1308 ] = 32'h2300932E;
  assign memory[ 1309 ] = 32'h9B2E932F;
  assign memory[ 1310 ] = 32'h00189C2F;
  assign memory[ 1311 ] = 32'hB0400021;
  assign memory[ 1312 ] = 32'h46C0BD70;
  assign memory[ 1313 ] = 32'hFFFFC000;
  assign memory[ 1314 ] = 32'hB08BB500;
  assign memory[ 1315 ] = 32'h91009001;
  assign memory[ 1316 ] = 32'h039B9B01;
  assign memory[ 1317 ] = 32'h00189900;
  assign memory[ 1318 ] = 32'hFBEEF000;
  assign memory[ 1319 ] = 32'h93070003;
  assign memory[ 1320 ] = 32'h681A4B2E;
  assign memory[ 1321 ] = 32'h429A9B07;
  assign memory[ 1322 ] = 32'h4B2CD903;
  assign memory[ 1323 ] = 32'h9309685B;
  assign memory[ 1324 ] = 32'h4B2AE050;
  assign memory[ 1325 ] = 32'h589A2298;
  assign memory[ 1326 ] = 32'h429A9B07;
  assign memory[ 1327 ] = 32'h4B27D804;
  assign memory[ 1328 ] = 32'h589B229C;
  assign memory[ 1329 ] = 32'hE0459309;
  assign memory[ 1330 ] = 32'h93082300;
  assign memory[ 1331 ] = 32'h4B23E03F;
  assign memory[ 1332 ] = 32'h00D29A08;
  assign memory[ 1333 ] = 32'h9B0758D2;
  assign memory[ 1334 ] = 32'hD835429A;
  assign memory[ 1335 ] = 32'h1C5A9B08;
  assign memory[ 1336 ] = 32'h00D24B1E;
  assign memory[ 1337 ] = 32'h9B0758D2;
  assign memory[ 1338 ] = 32'hD92D429A;
  assign memory[ 1339 ] = 32'h9A084B1B;
  assign memory[ 1340 ] = 32'h58D300D2;
  assign memory[ 1341 ] = 32'h9B089306;
  assign memory[ 1342 ] = 32'h4B181C5A;
  assign memory[ 1343 ] = 32'h58D300D2;
  assign memory[ 1344 ] = 32'h4A169305;
  assign memory[ 1345 ] = 32'h00DB9B08;
  assign memory[ 1346 ] = 32'h330418D3;
  assign memory[ 1347 ] = 32'h9304681B;
  assign memory[ 1348 ] = 32'h33019B08;
  assign memory[ 1349 ] = 32'h00DB4A11;
  assign memory[ 1350 ] = 32'h330418D3;
  assign memory[ 1351 ] = 32'h9303681B;
  assign memory[ 1352 ] = 32'h9B069A07;
  assign memory[ 1353 ] = 32'h99031AD3;
  assign memory[ 1354 ] = 32'h1A8A9A04;
  assign memory[ 1355 ] = 32'h0010435A;
  assign memory[ 1356 ] = 32'h9B069A05;
  assign memory[ 1357 ] = 32'h00191AD3;
  assign memory[ 1358 ] = 32'hFC28F000;
  assign memory[ 1359 ] = 32'h001A0003;
  assign memory[ 1360 ] = 32'h18D39B04;
  assign memory[ 1361 ] = 32'hE0059309;
  assign memory[ 1362 ] = 32'h33019B08;
  assign memory[ 1363 ] = 32'h9B089308;
  assign memory[ 1364 ] = 32'hDDBC2B12;
  assign memory[ 1365 ] = 32'h00189B09;
  assign memory[ 1366 ] = 32'hBD00B00B;
  assign memory[ 1367 ] = 32'h2000000C;
  assign memory[ 1368 ] = 32'h9001B082;
  assign memory[ 1369 ] = 32'h22204B13;
  assign memory[ 1370 ] = 32'h001A5C9B;
  assign memory[ 1371 ] = 32'h00924B11;
  assign memory[ 1372 ] = 32'h50D19901;
  assign memory[ 1373 ] = 32'h22204B0F;
  assign memory[ 1374 ] = 32'h33015C9B;
  assign memory[ 1375 ] = 32'h40134A0E;
  assign memory[ 1376 ] = 32'h3B01D504;
  assign memory[ 1377 ] = 32'h42522208;
  assign memory[ 1378 ] = 32'h33014313;
  assign memory[ 1379 ] = 32'h4B09B2D9;
  assign memory[ 1380 ] = 32'h54992220;
  assign memory[ 1381 ] = 32'h22214B07;
  assign memory[ 1382 ] = 32'h2B075C9B;
  assign memory[ 1383 ] = 32'h4B05D807;
  assign memory[ 1384 ] = 32'h5C9B2221;
  assign memory[ 1385 ] = 32'hB2D93301;
  assign memory[ 1386 ] = 32'h22214B02;
  assign memory[ 1387 ] = 32'h46C05499;
  assign memory[ 1388 ] = 32'h4770B002;
  assign memory[ 1389 ] = 32'h200000DC;
  assign memory[ 1390 ] = 32'h80000007;
  assign memory[ 1391 ] = 32'hB083B5F0;
  assign memory[ 1392 ] = 32'h22214B1E;
  assign memory[ 1393 ] = 32'h2B005C9B;
  assign memory[ 1394 ] = 32'h2300D101;
  assign memory[ 1395 ] = 32'h2300E033;
  assign memory[ 1396 ] = 32'h466B9301;
  assign memory[ 1397 ] = 32'h22003303;
  assign memory[ 1398 ] = 32'hE013701A;
  assign memory[ 1399 ] = 32'h3303466B;
  assign memory[ 1400 ] = 32'h4B16781A;
  assign memory[ 1401 ] = 32'h58D20092;
  assign memory[ 1402 ] = 32'h00119B01;
  assign memory[ 1403 ] = 32'hF7FE0018;
  assign memory[ 1404 ] = 32'h0003FDCB;
  assign memory[ 1405 ] = 32'h466B9301;
  assign memory[ 1406 ] = 32'h781A3303;
  assign memory[ 1407 ] = 32'h3303466B;
  assign memory[ 1408 ] = 32'h701A3201;
  assign memory[ 1409 ] = 32'h22214B0D;
  assign memory[ 1410 ] = 32'h466A5C9B;
  assign memory[ 1411 ] = 32'h78123203;
  assign memory[ 1412 ] = 32'hD3E3429A;
  assign memory[ 1413 ] = 32'h22214B09;
  assign memory[ 1414 ] = 32'h001E5C9B;
  assign memory[ 1415 ] = 32'h001F2300;
  assign memory[ 1416 ] = 32'h03BD0CB3;
  assign memory[ 1417 ] = 32'h03B4431D;
  assign memory[ 1418 ] = 32'h9B010022;
  assign memory[ 1419 ] = 32'h00180011;
  assign memory[ 1420 ] = 32'hFDBEF7FE;
  assign memory[ 1421 ] = 32'h00180003;
  assign memory[ 1422 ] = 32'hBDF0B003;
  assign memory[ 1423 ] = 32'h200000DC;
  assign memory[ 1424 ] = 32'hB08BB5F0;
  assign memory[ 1425 ] = 32'h20009005;
  assign memory[ 1426 ] = 32'hFF5AF7FE;
  assign memory[ 1427 ] = 32'h93090003;
  assign memory[ 1428 ] = 32'h93082300;
  assign memory[ 1429 ] = 32'h681B4B2D;
  assign memory[ 1430 ] = 32'h42934A2D;
  assign memory[ 1431 ] = 32'h9B09D04A;
  assign memory[ 1432 ] = 32'h23009300;
  assign memory[ 1433 ] = 32'h99009301;
  assign memory[ 1434 ] = 32'h000B9A01;
  assign memory[ 1435 ] = 32'h00100C9B;
  assign memory[ 1436 ] = 32'h431F0387;
  assign memory[ 1437 ] = 32'h039E000B;
  assign memory[ 1438 ] = 32'h4B240032;
  assign memory[ 1439 ] = 32'h9302681B;
  assign memory[ 1440 ] = 32'h93032300;
  assign memory[ 1441 ] = 32'h99039802;
  assign memory[ 1442 ] = 32'h0C9B0003;
  assign memory[ 1443 ] = 32'h03B5000E;
  assign memory[ 1444 ] = 32'h0003431D;
  assign memory[ 1445 ] = 32'h0023039C;
  assign memory[ 1446 ] = 32'h00100019;
  assign memory[ 1447 ] = 32'hFD7EF7FE;
  assign memory[ 1448 ] = 32'h93080003;
  assign memory[ 1449 ] = 32'h23809A08;
  assign memory[ 1450 ] = 32'h429A01DB;
  assign memory[ 1451 ] = 32'h4B19DD28;
  assign memory[ 1452 ] = 32'h9B05681A;
  assign memory[ 1453 ] = 32'h00180011;
  assign memory[ 1454 ] = 32'hFD70F7FE;
  assign memory[ 1455 ] = 32'h93070003;
  assign memory[ 1456 ] = 32'h9B079A08;
  assign memory[ 1457 ] = 32'h00180011;
  assign memory[ 1458 ] = 32'hFD72F7FE;
  assign memory[ 1459 ] = 32'h4B120002;
  assign memory[ 1460 ] = 32'h4B11601A;
  assign memory[ 1461 ] = 32'h0018681B;
  assign memory[ 1462 ] = 32'hFF42F7FF;
  assign memory[ 1463 ] = 32'hFF6EF7FF;
  assign memory[ 1464 ] = 32'h4B0E0002;
  assign memory[ 1465 ] = 32'h4B0B601A;
  assign memory[ 1466 ] = 32'h601A9A05;
  assign memory[ 1467 ] = 32'h9A094B07;
  assign memory[ 1468 ] = 32'hE005601A;
  assign memory[ 1469 ] = 32'h9A054B07;
  assign memory[ 1470 ] = 32'h4B04601A;
  assign memory[ 1471 ] = 32'h601A9A09;
  assign memory[ 1472 ] = 32'h681B4B06;
  assign memory[ 1473 ] = 32'hB00B0018;
  assign memory[ 1474 ] = 32'h46C0BDF0;
  assign memory[ 1475 ] = 32'h200000AC;
  assign memory[ 1476 ] = 32'h0012D687;
  assign memory[ 1477 ] = 32'h200000C4;
  assign memory[ 1478 ] = 32'h200000CC;
  assign memory[ 1479 ] = 32'h200000C8;
  assign memory[ 1480 ] = 32'h9001B082;
  assign memory[ 1481 ] = 32'h2B099B01;
  assign memory[ 1482 ] = 32'h2300D101;
  assign memory[ 1483 ] = 32'h9B01E001;
  assign memory[ 1484 ] = 32'h00183301;
  assign memory[ 1485 ] = 32'h4770B002;
  assign memory[ 1486 ] = 32'hB086B510;
  assign memory[ 1487 ] = 32'h0018466B;
  assign memory[ 1488 ] = 32'h001A2306;
  assign memory[ 1489 ] = 32'hF0002100;
  assign memory[ 1490 ] = 32'h2317FD81;
  assign memory[ 1491 ] = 32'h2205446B;
  assign memory[ 1492 ] = 32'h466B701A;
  assign memory[ 1493 ] = 32'hF7FF0018;
  assign memory[ 1494 ] = 32'h46C0FA4B;
  assign memory[ 1495 ] = 32'hFEA8F7FE;
  assign memory[ 1496 ] = 32'hD1FB1E03;
  assign memory[ 1497 ] = 32'hFF34F7FE;
  assign memory[ 1498 ] = 32'hF7FE46C0;
  assign memory[ 1499 ] = 32'h0003FD3D;
  assign memory[ 1500 ] = 32'h2301001A;
  assign memory[ 1501 ] = 32'hB2DB4053;
  assign memory[ 1502 ] = 32'hD1F62B00;
  assign memory[ 1503 ] = 32'hFD34F7FE;
  assign memory[ 1504 ] = 32'hD0131E03;
  assign memory[ 1505 ] = 32'hFD3CF7FE;
  assign memory[ 1506 ] = 32'h93020003;
  assign memory[ 1507 ] = 32'h22019B02;
  assign memory[ 1508 ] = 32'h230F401A;
  assign memory[ 1509 ] = 32'h1E51446B;
  assign memory[ 1510 ] = 32'h701A418A;
  assign memory[ 1511 ] = 32'h22029B02;
  assign memory[ 1512 ] = 32'h230E401A;
  assign memory[ 1513 ] = 32'h1E51446B;
  assign memory[ 1514 ] = 32'h701A418A;
  assign memory[ 1515 ] = 32'h446B230F;
  assign memory[ 1516 ] = 32'h2B00781B;
  assign memory[ 1517 ] = 32'h2317D00C;
  assign memory[ 1518 ] = 32'h781B446B;
  assign memory[ 1519 ] = 32'hD01C2B00;
  assign memory[ 1520 ] = 32'h446B2317;
  assign memory[ 1521 ] = 32'h446A2217;
  assign memory[ 1522 ] = 32'h3A017812;
  assign memory[ 1523 ] = 32'hE7C0701A;
  assign memory[ 1524 ] = 32'h446B230E;
  assign memory[ 1525 ] = 32'h2B00781B;
  assign memory[ 1526 ] = 32'h2317D0BB;
  assign memory[ 1527 ] = 32'h781C446B;
  assign memory[ 1528 ] = 32'h446B2317;
  assign memory[ 1529 ] = 32'h466A781B;
  assign memory[ 1530 ] = 32'h00185CD3;
  assign memory[ 1531 ] = 32'hFF98F7FF;
  assign memory[ 1532 ] = 32'hB2DA0003;
  assign memory[ 1533 ] = 32'h551A466B;
  assign memory[ 1534 ] = 32'h46C0E7AB;
  assign memory[ 1535 ] = 32'h795B466B;
  assign memory[ 1536 ] = 32'h4B15001A;
  assign memory[ 1537 ] = 32'h466B435A;
  assign memory[ 1538 ] = 32'h0019791B;
  assign memory[ 1539 ] = 32'h434B4B13;
  assign memory[ 1540 ] = 32'h466B18D2;
  assign memory[ 1541 ] = 32'h001978DB;
  assign memory[ 1542 ] = 32'h009B23FA;
  assign memory[ 1543 ] = 32'h18D2434B;
  assign memory[ 1544 ] = 32'h789B466B;
  assign memory[ 1545 ] = 32'h23640019;
  assign memory[ 1546 ] = 32'h18D2434B;
  assign memory[ 1547 ] = 32'h785B466B;
  assign memory[ 1548 ] = 32'h000B0019;
  assign memory[ 1549 ] = 32'h185B009B;
  assign memory[ 1550 ] = 32'h18D3005B;
  assign memory[ 1551 ] = 32'h7812466A;
  assign memory[ 1552 ] = 32'h9304189B;
  assign memory[ 1553 ] = 32'h2B009B04;
  assign memory[ 1554 ] = 32'h4B05D101;
  assign memory[ 1555 ] = 32'h9B049304;
  assign memory[ 1556 ] = 32'hB0060018;
  assign memory[ 1557 ] = 32'h46C0BD10;
  assign memory[ 1558 ] = 32'h000186A0;
  assign memory[ 1559 ] = 32'h00002710;
  assign memory[ 1560 ] = 32'h00018BCD;
  assign memory[ 1561 ] = 32'hB084B510;
  assign memory[ 1562 ] = 32'h2200466B;
  assign memory[ 1563 ] = 32'h230F601A;
  assign memory[ 1564 ] = 32'h2203446B;
  assign memory[ 1565 ] = 32'h466B701A;
  assign memory[ 1566 ] = 32'hF7FF0018;
  assign memory[ 1567 ] = 32'h46C0FA27;
  assign memory[ 1568 ] = 32'hFE16F7FE;
  assign memory[ 1569 ] = 32'hD1FB1E03;
  assign memory[ 1570 ] = 32'hFEA2F7FE;
  assign memory[ 1571 ] = 32'hF7FE46C0;
  assign memory[ 1572 ] = 32'h0003FCAB;
  assign memory[ 1573 ] = 32'h2301001A;
  assign memory[ 1574 ] = 32'hB2DB4053;
  assign memory[ 1575 ] = 32'hD1F62B00;
  assign memory[ 1576 ] = 32'hFCA2F7FE;
  assign memory[ 1577 ] = 32'hD0131E03;
  assign memory[ 1578 ] = 32'hFCAAF7FE;
  assign memory[ 1579 ] = 32'h93020003;
  assign memory[ 1580 ] = 32'h22019B02;
  assign memory[ 1581 ] = 32'h230E401A;
  assign memory[ 1582 ] = 32'h1E51446B;
  assign memory[ 1583 ] = 32'h701A418A;
  assign memory[ 1584 ] = 32'h22029B02;
  assign memory[ 1585 ] = 32'h230D401A;
  assign memory[ 1586 ] = 32'h1E51446B;
  assign memory[ 1587 ] = 32'h701A418A;
  assign memory[ 1588 ] = 32'h446B230E;
  assign memory[ 1589 ] = 32'h2B00781B;
  assign memory[ 1590 ] = 32'h230FD00C;
  assign memory[ 1591 ] = 32'h781B446B;
  assign memory[ 1592 ] = 32'hD01C2B00;
  assign memory[ 1593 ] = 32'h446B230F;
  assign memory[ 1594 ] = 32'h446A220F;
  assign memory[ 1595 ] = 32'h3A017812;
  assign memory[ 1596 ] = 32'hE7C0701A;
  assign memory[ 1597 ] = 32'h446B230D;
  assign memory[ 1598 ] = 32'h2B00781B;
  assign memory[ 1599 ] = 32'h230FD0BB;
  assign memory[ 1600 ] = 32'h781C446B;
  assign memory[ 1601 ] = 32'h446B230F;
  assign memory[ 1602 ] = 32'h466A781B;
  assign memory[ 1603 ] = 32'h00185CD3;
  assign memory[ 1604 ] = 32'hFF06F7FF;
  assign memory[ 1605 ] = 32'hB2DA0003;
  assign memory[ 1606 ] = 32'h551A466B;
  assign memory[ 1607 ] = 32'h46C0E7AB;
  assign memory[ 1608 ] = 32'h78DB466B;
  assign memory[ 1609 ] = 32'h23FA001A;
  assign memory[ 1610 ] = 32'h435A009B;
  assign memory[ 1611 ] = 32'h789B466B;
  assign memory[ 1612 ] = 32'h23640019;
  assign memory[ 1613 ] = 32'h18D2434B;
  assign memory[ 1614 ] = 32'h785B466B;
  assign memory[ 1615 ] = 32'h000B0019;
  assign memory[ 1616 ] = 32'h185B009B;
  assign memory[ 1617 ] = 32'h18D3005B;
  assign memory[ 1618 ] = 32'h7812466A;
  assign memory[ 1619 ] = 32'h9301189B;
  assign memory[ 1620 ] = 32'h00189B01;
  assign memory[ 1621 ] = 32'hBD10B004;
  assign memory[ 1622 ] = 32'hB09BB5F0;
  assign memory[ 1623 ] = 32'h021B2380;
  assign memory[ 1624 ] = 32'hF7FE0018;
  assign memory[ 1625 ] = 32'hAB04FDBB;
  assign memory[ 1626 ] = 32'h23060018;
  assign memory[ 1627 ] = 32'h2100001A;
  assign memory[ 1628 ] = 32'hFC6CF000;
  assign memory[ 1629 ] = 32'hFE34F7FE;
  assign memory[ 1630 ] = 32'hF7FE2077;
  assign memory[ 1631 ] = 32'hF7FFFC71;
  assign memory[ 1632 ] = 32'h4BB8FA05;
  assign memory[ 1633 ] = 32'hF7FF0018;
  assign memory[ 1634 ] = 32'h2300FAB1;
  assign memory[ 1635 ] = 32'h4BB69318;
  assign memory[ 1636 ] = 32'h23009317;
  assign memory[ 1637 ] = 32'h23009316;
  assign memory[ 1638 ] = 32'hAB049313;
  assign memory[ 1639 ] = 32'h00192206;
  assign memory[ 1640 ] = 32'hF7FF2004;
  assign memory[ 1641 ] = 32'hAB04FA0B;
  assign memory[ 1642 ] = 32'h041A789B;
  assign memory[ 1643 ] = 32'h785BAB04;
  assign memory[ 1644 ] = 32'h18D3021B;
  assign memory[ 1645 ] = 32'h7812AA04;
  assign memory[ 1646 ] = 32'h9312189B;
  assign memory[ 1647 ] = 32'h795BAB04;
  assign memory[ 1648 ] = 32'hAB04041A;
  assign memory[ 1649 ] = 32'h021B791B;
  assign memory[ 1650 ] = 32'hAA0418D3;
  assign memory[ 1651 ] = 32'h189B78D2;
  assign memory[ 1652 ] = 32'h4AA49311;
  assign memory[ 1653 ] = 32'h00119B11;
  assign memory[ 1654 ] = 32'hF7FF0018;
  assign memory[ 1655 ] = 32'h0002FB19;
  assign memory[ 1656 ] = 32'h920E000B;
  assign memory[ 1657 ] = 32'h4A9F930F;
  assign memory[ 1658 ] = 32'h00119B12;
  assign memory[ 1659 ] = 32'hF7FF0018;
  assign memory[ 1660 ] = 32'h0002FB7F;
  assign memory[ 1661 ] = 32'h920C000B;
  assign memory[ 1662 ] = 32'h9B0C930D;
  assign memory[ 1663 ] = 32'h00119A17;
  assign memory[ 1664 ] = 32'hF7FF0018;
  assign memory[ 1665 ] = 32'h0003FD41;
  assign memory[ 1666 ] = 32'h9B169316;
  assign memory[ 1667 ] = 32'h23009300;
  assign memory[ 1668 ] = 32'h99009301;
  assign memory[ 1669 ] = 32'h000B9A01;
  assign memory[ 1670 ] = 32'h00100C9B;
  assign memory[ 1671 ] = 32'h431D0385;
  assign memory[ 1672 ] = 32'h039C000B;
  assign memory[ 1673 ] = 32'h00180023;
  assign memory[ 1674 ] = 32'hFE0AF7FF;
  assign memory[ 1675 ] = 32'h93130003;
  assign memory[ 1676 ] = 32'h4A8E9B16;
  assign memory[ 1677 ] = 32'hD9014293;
  assign memory[ 1678 ] = 32'h93164B8C;
  assign memory[ 1679 ] = 32'hAA042357;
  assign memory[ 1680 ] = 32'h44634694;
  assign memory[ 1681 ] = 32'h701A2200;
  assign memory[ 1682 ] = 32'hAA042356;
  assign memory[ 1683 ] = 32'h44634694;
  assign memory[ 1684 ] = 32'h701A2200;
  assign memory[ 1685 ] = 32'hAA042355;
  assign memory[ 1686 ] = 32'h44634694;
  assign memory[ 1687 ] = 32'h701A2200;
  assign memory[ 1688 ] = 32'hFBC2F7FE;
  assign memory[ 1689 ] = 32'hD0211E03;
  assign memory[ 1690 ] = 32'hFBCAF7FE;
  assign memory[ 1691 ] = 32'h930B0003;
  assign memory[ 1692 ] = 32'h22019B0B;
  assign memory[ 1693 ] = 32'h2357401A;
  assign memory[ 1694 ] = 32'h468CA904;
  assign memory[ 1695 ] = 32'h1E514463;
  assign memory[ 1696 ] = 32'h701A418A;
  assign memory[ 1697 ] = 32'h22029B0B;
  assign memory[ 1698 ] = 32'h2356401A;
  assign memory[ 1699 ] = 32'h468CA904;
  assign memory[ 1700 ] = 32'h1E514463;
  assign memory[ 1701 ] = 32'h701A418A;
  assign memory[ 1702 ] = 32'h22049B0B;
  assign memory[ 1703 ] = 32'h2355401A;
  assign memory[ 1704 ] = 32'h468CA904;
  assign memory[ 1705 ] = 32'h1E514463;
  assign memory[ 1706 ] = 32'h701A418A;
  assign memory[ 1707 ] = 32'hAA042357;
  assign memory[ 1708 ] = 32'h44634694;
  assign memory[ 1709 ] = 32'h2B00781B;
  assign memory[ 1710 ] = 32'h9B18D017;
  assign memory[ 1711 ] = 32'hD0082B01;
  assign memory[ 1712 ] = 32'h2B02D304;
  assign memory[ 1713 ] = 32'h2B03D008;
  assign memory[ 1714 ] = 32'hE00BD009;
  assign memory[ 1715 ] = 32'h93182301;
  assign memory[ 1716 ] = 32'h2302E00B;
  assign memory[ 1717 ] = 32'hE0089318;
  assign memory[ 1718 ] = 32'h93182303;
  assign memory[ 1719 ] = 32'h2300E005;
  assign memory[ 1720 ] = 32'hE0029318;
  assign memory[ 1721 ] = 32'h93182300;
  assign memory[ 1722 ] = 32'h235646C0;
  assign memory[ 1723 ] = 32'h4694AA04;
  assign memory[ 1724 ] = 32'h781B4463;
  assign memory[ 1725 ] = 32'hD0022B00;
  assign memory[ 1726 ] = 32'h22004B5D;
  assign memory[ 1727 ] = 32'h2355601A;
  assign memory[ 1728 ] = 32'h4694AA04;
  assign memory[ 1729 ] = 32'h781B4463;
  assign memory[ 1730 ] = 32'hD1002B00;
  assign memory[ 1731 ] = 32'h9B18E081;
  assign memory[ 1732 ] = 32'hD1032B00;
  assign memory[ 1733 ] = 32'hFE10F7FF;
  assign memory[ 1734 ] = 32'h93170003;
  assign memory[ 1735 ] = 32'h2B019B18;
  assign memory[ 1736 ] = 32'hE076D000;
  assign memory[ 1737 ] = 32'hFE9EF7FF;
  assign memory[ 1738 ] = 32'h930A0003;
  assign memory[ 1739 ] = 32'h685A4B51;
  assign memory[ 1740 ] = 32'h429A9B0A;
  assign memory[ 1741 ] = 32'h4B4FD803;
  assign memory[ 1742 ] = 32'h9315681B;
  assign memory[ 1743 ] = 32'h4B4DE054;
  assign memory[ 1744 ] = 32'h589A229C;
  assign memory[ 1745 ] = 32'h429A9B0A;
  assign memory[ 1746 ] = 32'h4B4AD904;
  assign memory[ 1747 ] = 32'h589B2298;
  assign memory[ 1748 ] = 32'hE0499315;
  assign memory[ 1749 ] = 32'h93142300;
  assign memory[ 1750 ] = 32'h4A46E043;
  assign memory[ 1751 ] = 32'h00DB9B14;
  assign memory[ 1752 ] = 32'h330418D3;
  assign memory[ 1753 ] = 32'h9B0A681A;
  assign memory[ 1754 ] = 32'hD937429A;
  assign memory[ 1755 ] = 32'h33019B14;
  assign memory[ 1756 ] = 32'h00DB4A40;
  assign memory[ 1757 ] = 32'h330418D3;
  assign memory[ 1758 ] = 32'h9B0A681A;
  assign memory[ 1759 ] = 32'hD82D429A;
  assign memory[ 1760 ] = 32'h9A144B3C;
  assign memory[ 1761 ] = 32'h58D300D2;
  assign memory[ 1762 ] = 32'h9B149309;
  assign memory[ 1763 ] = 32'h4B391C5A;
  assign memory[ 1764 ] = 32'h58D300D2;
  assign memory[ 1765 ] = 32'h4A379308;
  assign memory[ 1766 ] = 32'h00DB9B14;
  assign memory[ 1767 ] = 32'h330418D3;
  assign memory[ 1768 ] = 32'h9307681B;
  assign memory[ 1769 ] = 32'h33019B14;
  assign memory[ 1770 ] = 32'h00DB4A32;
  assign memory[ 1771 ] = 32'h330418D3;
  assign memory[ 1772 ] = 32'h9306681B;
  assign memory[ 1773 ] = 32'h9B079A0A;
  assign memory[ 1774 ] = 32'h99081AD3;
  assign memory[ 1775 ] = 32'h1A8A9A09;
  assign memory[ 1776 ] = 32'h0010435A;
  assign memory[ 1777 ] = 32'h9B079A06;
  assign memory[ 1778 ] = 32'h00191AD3;
  assign memory[ 1779 ] = 32'hF8DEF000;
  assign memory[ 1780 ] = 32'h001A0003;
  assign memory[ 1781 ] = 32'h18D39B09;
  assign memory[ 1782 ] = 32'hE0059315;
  assign memory[ 1783 ] = 32'h33019B14;
  assign memory[ 1784 ] = 32'h9B149314;
  assign memory[ 1785 ] = 32'hDDB82B12;
  assign memory[ 1786 ] = 32'h0C9B9B0C;
  assign memory[ 1787 ] = 32'h03979A0D;
  assign memory[ 1788 ] = 32'h9B0C431F;
  assign memory[ 1789 ] = 32'h9B15039E;
  assign memory[ 1790 ] = 32'h17DB9302;
  assign memory[ 1791 ] = 32'h9A029303;
  assign memory[ 1792 ] = 32'h00309B03;
  assign memory[ 1793 ] = 32'hF0000039;
  assign memory[ 1794 ] = 32'h0002F9AD;
  assign memory[ 1795 ] = 32'h0013000B;
  assign memory[ 1796 ] = 32'h9B189317;
  assign memory[ 1797 ] = 32'hD00A2B01;
  assign memory[ 1798 ] = 32'h2B02D304;
  assign memory[ 1799 ] = 32'h2B03D00C;
  assign memory[ 1800 ] = 32'hE016D012;
  assign memory[ 1801 ] = 32'h00189B0C;
  assign memory[ 1802 ] = 32'hFD82F7FE;
  assign memory[ 1803 ] = 32'h9B16E011;
  assign memory[ 1804 ] = 32'hF7FE0018;
  assign memory[ 1805 ] = 32'hE00CFE1D;
  assign memory[ 1806 ] = 32'hF7FE2000;
  assign memory[ 1807 ] = 32'h0003FC61;
  assign memory[ 1808 ] = 32'hF7FE0018;
  assign memory[ 1809 ] = 32'hE004FEAD;
  assign memory[ 1810 ] = 32'h00189B13;
  assign memory[ 1811 ] = 32'hFF44F7FE;
  assign memory[ 1812 ] = 32'h46C046C0;
  assign memory[ 1813 ] = 32'hFC2CF7FE;
  assign memory[ 1814 ] = 32'hD1FB1E03;
  assign memory[ 1815 ] = 32'hFCB8F7FE;
  assign memory[ 1816 ] = 32'h46C0E69B;
  assign memory[ 1817 ] = 32'h20000100;
  assign memory[ 1818 ] = 32'h00018BCD;
  assign memory[ 1819 ] = 32'h0000270F;
  assign memory[ 1820 ] = 32'h200000C0;
  assign memory[ 1821 ] = 32'h2000000C;
  assign memory[ 1822 ] = 32'h08432200;
  assign memory[ 1823 ] = 32'hD374428B;
  assign memory[ 1824 ] = 32'h428B0903;
  assign memory[ 1825 ] = 32'h0A03D35F;
  assign memory[ 1826 ] = 32'hD344428B;
  assign memory[ 1827 ] = 32'h428B0B03;
  assign memory[ 1828 ] = 32'h0C03D328;
  assign memory[ 1829 ] = 32'hD30D428B;
  assign memory[ 1830 ] = 32'h020922FF;
  assign memory[ 1831 ] = 32'h0C03BA12;
  assign memory[ 1832 ] = 32'hD302428B;
  assign memory[ 1833 ] = 32'h02091212;
  assign memory[ 1834 ] = 32'h0B03D065;
  assign memory[ 1835 ] = 32'hD319428B;
  assign memory[ 1836 ] = 32'h0A09E000;
  assign memory[ 1837 ] = 32'h428B0BC3;
  assign memory[ 1838 ] = 32'h03CBD301;
  assign memory[ 1839 ] = 32'h41521AC0;
  assign memory[ 1840 ] = 32'h428B0B83;
  assign memory[ 1841 ] = 32'h038BD301;
  assign memory[ 1842 ] = 32'h41521AC0;
  assign memory[ 1843 ] = 32'h428B0B43;
  assign memory[ 1844 ] = 32'h034BD301;
  assign memory[ 1845 ] = 32'h41521AC0;
  assign memory[ 1846 ] = 32'h428B0B03;
  assign memory[ 1847 ] = 32'h030BD301;
  assign memory[ 1848 ] = 32'h41521AC0;
  assign memory[ 1849 ] = 32'h428B0AC3;
  assign memory[ 1850 ] = 32'h02CBD301;
  assign memory[ 1851 ] = 32'h41521AC0;
  assign memory[ 1852 ] = 32'h428B0A83;
  assign memory[ 1853 ] = 32'h028BD301;
  assign memory[ 1854 ] = 32'h41521AC0;
  assign memory[ 1855 ] = 32'h428B0A43;
  assign memory[ 1856 ] = 32'h024BD301;
  assign memory[ 1857 ] = 32'h41521AC0;
  assign memory[ 1858 ] = 32'h428B0A03;
  assign memory[ 1859 ] = 32'h020BD301;
  assign memory[ 1860 ] = 32'h41521AC0;
  assign memory[ 1861 ] = 32'h09C3D2CD;
  assign memory[ 1862 ] = 32'hD301428B;
  assign memory[ 1863 ] = 32'h1AC001CB;
  assign memory[ 1864 ] = 32'h09834152;
  assign memory[ 1865 ] = 32'hD301428B;
  assign memory[ 1866 ] = 32'h1AC0018B;
  assign memory[ 1867 ] = 32'h09434152;
  assign memory[ 1868 ] = 32'hD301428B;
  assign memory[ 1869 ] = 32'h1AC0014B;
  assign memory[ 1870 ] = 32'h09034152;
  assign memory[ 1871 ] = 32'hD301428B;
  assign memory[ 1872 ] = 32'h1AC0010B;
  assign memory[ 1873 ] = 32'h08C34152;
  assign memory[ 1874 ] = 32'hD301428B;
  assign memory[ 1875 ] = 32'h1AC000CB;
  assign memory[ 1876 ] = 32'h08834152;
  assign memory[ 1877 ] = 32'hD301428B;
  assign memory[ 1878 ] = 32'h1AC0008B;
  assign memory[ 1879 ] = 32'h08434152;
  assign memory[ 1880 ] = 32'hD301428B;
  assign memory[ 1881 ] = 32'h1AC0004B;
  assign memory[ 1882 ] = 32'h1A414152;
  assign memory[ 1883 ] = 32'h4601D200;
  assign memory[ 1884 ] = 32'h46104152;
  assign memory[ 1885 ] = 32'hE7FF4770;
  assign memory[ 1886 ] = 32'h2000B501;
  assign memory[ 1887 ] = 32'hF8F0F000;
  assign memory[ 1888 ] = 32'h46C0BD02;
  assign memory[ 1889 ] = 32'hD0F72900;
  assign memory[ 1890 ] = 32'h4770E776;
  assign memory[ 1891 ] = 32'h430B4603;
  assign memory[ 1892 ] = 32'h2200D47F;
  assign memory[ 1893 ] = 32'h428B0843;
  assign memory[ 1894 ] = 32'h0903D374;
  assign memory[ 1895 ] = 32'hD35F428B;
  assign memory[ 1896 ] = 32'h428B0A03;
  assign memory[ 1897 ] = 32'h0B03D344;
  assign memory[ 1898 ] = 32'hD328428B;
  assign memory[ 1899 ] = 32'h428B0C03;
  assign memory[ 1900 ] = 32'h22FFD30D;
  assign memory[ 1901 ] = 32'hBA120209;
  assign memory[ 1902 ] = 32'h428B0C03;
  assign memory[ 1903 ] = 32'h1212D302;
  assign memory[ 1904 ] = 32'hD0650209;
  assign memory[ 1905 ] = 32'h428B0B03;
  assign memory[ 1906 ] = 32'hE000D319;
  assign memory[ 1907 ] = 32'h0BC30A09;
  assign memory[ 1908 ] = 32'hD301428B;
  assign memory[ 1909 ] = 32'h1AC003CB;
  assign memory[ 1910 ] = 32'h0B834152;
  assign memory[ 1911 ] = 32'hD301428B;
  assign memory[ 1912 ] = 32'h1AC0038B;
  assign memory[ 1913 ] = 32'h0B434152;
  assign memory[ 1914 ] = 32'hD301428B;
  assign memory[ 1915 ] = 32'h1AC0034B;
  assign memory[ 1916 ] = 32'h0B034152;
  assign memory[ 1917 ] = 32'hD301428B;
  assign memory[ 1918 ] = 32'h1AC0030B;
  assign memory[ 1919 ] = 32'h0AC34152;
  assign memory[ 1920 ] = 32'hD301428B;
  assign memory[ 1921 ] = 32'h1AC002CB;
  assign memory[ 1922 ] = 32'h0A834152;
  assign memory[ 1923 ] = 32'hD301428B;
  assign memory[ 1924 ] = 32'h1AC0028B;
  assign memory[ 1925 ] = 32'h0A434152;
  assign memory[ 1926 ] = 32'hD301428B;
  assign memory[ 1927 ] = 32'h1AC0024B;
  assign memory[ 1928 ] = 32'h0A034152;
  assign memory[ 1929 ] = 32'hD301428B;
  assign memory[ 1930 ] = 32'h1AC0020B;
  assign memory[ 1931 ] = 32'hD2CD4152;
  assign memory[ 1932 ] = 32'h428B09C3;
  assign memory[ 1933 ] = 32'h01CBD301;
  assign memory[ 1934 ] = 32'h41521AC0;
  assign memory[ 1935 ] = 32'h428B0983;
  assign memory[ 1936 ] = 32'h018BD301;
  assign memory[ 1937 ] = 32'h41521AC0;
  assign memory[ 1938 ] = 32'h428B0943;
  assign memory[ 1939 ] = 32'h014BD301;
  assign memory[ 1940 ] = 32'h41521AC0;
  assign memory[ 1941 ] = 32'h428B0903;
  assign memory[ 1942 ] = 32'h010BD301;
  assign memory[ 1943 ] = 32'h41521AC0;
  assign memory[ 1944 ] = 32'h428B08C3;
  assign memory[ 1945 ] = 32'h00CBD301;
  assign memory[ 1946 ] = 32'h41521AC0;
  assign memory[ 1947 ] = 32'h428B0883;
  assign memory[ 1948 ] = 32'h008BD301;
  assign memory[ 1949 ] = 32'h41521AC0;
  assign memory[ 1950 ] = 32'h428B0843;
  assign memory[ 1951 ] = 32'h004BD301;
  assign memory[ 1952 ] = 32'h41521AC0;
  assign memory[ 1953 ] = 32'hD2001A41;
  assign memory[ 1954 ] = 32'h41524601;
  assign memory[ 1955 ] = 32'h47704610;
  assign memory[ 1956 ] = 32'h0FCAE05D;
  assign memory[ 1957 ] = 32'h4249D000;
  assign memory[ 1958 ] = 32'hD3001003;
  assign memory[ 1959 ] = 32'h40534240;
  assign memory[ 1960 ] = 32'h469C2200;
  assign memory[ 1961 ] = 32'h428B0903;
  assign memory[ 1962 ] = 32'h0A03D32D;
  assign memory[ 1963 ] = 32'hD312428B;
  assign memory[ 1964 ] = 32'h018922FC;
  assign memory[ 1965 ] = 32'h0A03BA12;
  assign memory[ 1966 ] = 32'hD30C428B;
  assign memory[ 1967 ] = 32'h11920189;
  assign memory[ 1968 ] = 32'hD308428B;
  assign memory[ 1969 ] = 32'h11920189;
  assign memory[ 1970 ] = 32'hD304428B;
  assign memory[ 1971 ] = 32'hD03A0189;
  assign memory[ 1972 ] = 32'hE0001192;
  assign memory[ 1973 ] = 32'h09C30989;
  assign memory[ 1974 ] = 32'hD301428B;
  assign memory[ 1975 ] = 32'h1AC001CB;
  assign memory[ 1976 ] = 32'h09834152;
  assign memory[ 1977 ] = 32'hD301428B;
  assign memory[ 1978 ] = 32'h1AC0018B;
  assign memory[ 1979 ] = 32'h09434152;
  assign memory[ 1980 ] = 32'hD301428B;
  assign memory[ 1981 ] = 32'h1AC0014B;
  assign memory[ 1982 ] = 32'h09034152;
  assign memory[ 1983 ] = 32'hD301428B;
  assign memory[ 1984 ] = 32'h1AC0010B;
  assign memory[ 1985 ] = 32'h08C34152;
  assign memory[ 1986 ] = 32'hD301428B;
  assign memory[ 1987 ] = 32'h1AC000CB;
  assign memory[ 1988 ] = 32'h08834152;
  assign memory[ 1989 ] = 32'hD301428B;
  assign memory[ 1990 ] = 32'h1AC0008B;
  assign memory[ 1991 ] = 32'hD2D94152;
  assign memory[ 1992 ] = 32'h428B0843;
  assign memory[ 1993 ] = 32'h004BD301;
  assign memory[ 1994 ] = 32'h41521AC0;
  assign memory[ 1995 ] = 32'hD2001A41;
  assign memory[ 1996 ] = 32'h46634601;
  assign memory[ 1997 ] = 32'h105B4152;
  assign memory[ 1998 ] = 32'hD3014610;
  assign memory[ 1999 ] = 32'h2B004240;
  assign memory[ 2000 ] = 32'h4249D500;
  assign memory[ 2001 ] = 32'h46634770;
  assign memory[ 2002 ] = 32'hD300105B;
  assign memory[ 2003 ] = 32'hB5014240;
  assign memory[ 2004 ] = 32'hF0002000;
  assign memory[ 2005 ] = 32'hBD02F805;
  assign memory[ 2006 ] = 32'hD0F82900;
  assign memory[ 2007 ] = 32'h4770E716;
  assign memory[ 2008 ] = 32'h46C04770;
  assign memory[ 2009 ] = 32'hD1152B00;
  assign memory[ 2010 ] = 32'hD1132A00;
  assign memory[ 2011 ] = 32'hDB062900;
  assign memory[ 2012 ] = 32'h2800DC01;
  assign memory[ 2013 ] = 32'h2000D006;
  assign memory[ 2014 ] = 32'h084143C0;
  assign memory[ 2015 ] = 32'h2180E002;
  assign memory[ 2016 ] = 32'h20000609;
  assign memory[ 2017 ] = 32'h4802B407;
  assign memory[ 2018 ] = 32'h1840A101;
  assign memory[ 2019 ] = 32'hBD039002;
  assign memory[ 2020 ] = 32'hFFFFFFD1;
  assign memory[ 2021 ] = 32'h4668B403;
  assign memory[ 2022 ] = 32'h9802B501;
  assign memory[ 2023 ] = 32'hF832F000;
  assign memory[ 2024 ] = 32'h469E9B01;
  assign memory[ 2025 ] = 32'hBC0CB002;
  assign memory[ 2026 ] = 32'h46C04770;
  assign memory[ 2027 ] = 32'h464FB5F0;
  assign memory[ 2028 ] = 32'hB4C04646;
  assign memory[ 2029 ] = 32'h0C360416;
  assign memory[ 2030 ] = 32'h00334699;
  assign memory[ 2031 ] = 32'h0C2C0405;
  assign memory[ 2032 ] = 32'h0C150C07;
  assign memory[ 2033 ] = 32'h437E4363;
  assign memory[ 2034 ] = 32'h4365436F;
  assign memory[ 2035 ] = 32'h19AD0C1C;
  assign memory[ 2036 ] = 32'h469C1964;
  assign memory[ 2037 ] = 32'hD90342A6;
  assign memory[ 2038 ] = 32'h025B2380;
  assign memory[ 2039 ] = 32'h44474698;
  assign memory[ 2040 ] = 32'h0C254663;
  assign memory[ 2041 ] = 32'h041D19EF;
  assign memory[ 2042 ] = 32'h434A464B;
  assign memory[ 2043 ] = 32'h0C2D4343;
  assign memory[ 2044 ] = 32'h19640424;
  assign memory[ 2045 ] = 32'h19C91899;
  assign memory[ 2046 ] = 32'hBC0C0020;
  assign memory[ 2047 ] = 32'h46994690;
  assign memory[ 2048 ] = 32'h46C0BDF0;
  assign memory[ 2049 ] = 32'hB083B5F0;
  assign memory[ 2050 ] = 32'h001F0016;
  assign memory[ 2051 ] = 32'h91019000;
  assign memory[ 2052 ] = 32'hF814F000;
  assign memory[ 2053 ] = 32'h000D0004;
  assign memory[ 2054 ] = 32'h000B0002;
  assign memory[ 2055 ] = 32'h00390030;
  assign memory[ 2056 ] = 32'hFFC4F7FF;
  assign memory[ 2057 ] = 32'h9B019A00;
  assign memory[ 2058 ] = 32'h418B1A12;
  assign memory[ 2059 ] = 32'h00209908;
  assign memory[ 2060 ] = 32'h604B600A;
  assign memory[ 2061 ] = 32'hB0030029;
  assign memory[ 2062 ] = 32'h46C0BDF0;
  assign memory[ 2063 ] = 32'h4644B5F0;
  assign memory[ 2064 ] = 32'h4656465F;
  assign memory[ 2065 ] = 32'hB4F0464D;
  assign memory[ 2066 ] = 32'hB083001C;
  assign memory[ 2067 ] = 32'hDA002900;
  assign memory[ 2068 ] = 32'h000FE092;
  assign memory[ 2069 ] = 32'h00062100;
  assign memory[ 2070 ] = 32'h0010468A;
  assign memory[ 2071 ] = 32'h2C000019;
  assign memory[ 2072 ] = 32'hE080DA00;
  assign memory[ 2073 ] = 32'h003D0034;
  assign memory[ 2074 ] = 32'h46884681;
  assign memory[ 2075 ] = 32'hD86942B9;
  assign memory[ 2076 ] = 32'h4641D066;
  assign memory[ 2077 ] = 32'hF0004648;
  assign memory[ 2078 ] = 32'h4683F8BF;
  assign memory[ 2079 ] = 32'h00300039;
  assign memory[ 2080 ] = 32'hF8BAF000;
  assign memory[ 2081 ] = 32'h1A1B465B;
  assign memory[ 2082 ] = 32'h3B20469C;
  assign memory[ 2083 ] = 32'hD500469B;
  assign memory[ 2084 ] = 32'h4649E086;
  assign memory[ 2085 ] = 32'h40814658;
  assign memory[ 2086 ] = 32'h4649000B;
  assign memory[ 2087 ] = 32'h40814660;
  assign memory[ 2088 ] = 32'h42BB000A;
  assign memory[ 2089 ] = 32'hE071D900;
  assign memory[ 2090 ] = 32'h0034D06D;
  assign memory[ 2091 ] = 32'h4659003D;
  assign memory[ 2092 ] = 32'h419D1AA4;
  assign memory[ 2093 ] = 32'hDA002900;
  assign memory[ 2094 ] = 32'h2100E089;
  assign memory[ 2095 ] = 32'h26012000;
  assign memory[ 2096 ] = 32'h91019000;
  assign memory[ 2097 ] = 32'h408E4659;
  assign memory[ 2098 ] = 32'h46619601;
  assign memory[ 2099 ] = 32'h408E2601;
  assign memory[ 2100 ] = 32'h96004661;
  assign memory[ 2101 ] = 32'hD0602900;
  assign memory[ 2102 ] = 32'h085607D9;
  assign memory[ 2103 ] = 32'h085F430E;
  assign memory[ 2104 ] = 32'h22014661;
  assign memory[ 2105 ] = 32'hE00C2300;
  assign memory[ 2106 ] = 32'hD10142AF;
  assign memory[ 2107 ] = 32'hD80A42A6;
  assign memory[ 2108 ] = 32'h41BD1BA4;
  assign memory[ 2109 ] = 32'h416D1924;
  assign memory[ 2110 ] = 32'h18A43901;
  assign memory[ 2111 ] = 32'h2900415D;
  assign memory[ 2112 ] = 32'h42AFD006;
  assign memory[ 2113 ] = 32'h3901D9F0;
  assign memory[ 2114 ] = 32'h416D1924;
  assign memory[ 2115 ] = 32'hD1F82900;
  assign memory[ 2116 ] = 32'h9800465B;
  assign memory[ 2117 ] = 32'h19009901;
  assign memory[ 2118 ] = 32'h2B004169;
  assign memory[ 2119 ] = 32'h002EDB4C;
  assign memory[ 2120 ] = 32'h466340DE;
  assign memory[ 2121 ] = 32'h40DC002C;
  assign memory[ 2122 ] = 32'h2B00465B;
  assign memory[ 2123 ] = 32'h0034DB5A;
  assign memory[ 2124 ] = 32'h0023409C;
  assign memory[ 2125 ] = 32'h40A64664;
  assign memory[ 2126 ] = 32'h1A800032;
  assign memory[ 2127 ] = 32'hE0034199;
  assign memory[ 2128 ] = 32'hD99642B0;
  assign memory[ 2129 ] = 32'h21002000;
  assign memory[ 2130 ] = 32'h2B004653;
  assign memory[ 2131 ] = 32'h0003D004;
  assign memory[ 2132 ] = 32'h2100000C;
  assign memory[ 2133 ] = 32'h41A14258;
  assign memory[ 2134 ] = 32'hBC3CB003;
  assign memory[ 2135 ] = 32'h46994690;
  assign memory[ 2136 ] = 32'h46AB46A2;
  assign memory[ 2137 ] = 32'h4653BDF0;
  assign memory[ 2138 ] = 32'h000C43DB;
  assign memory[ 2139 ] = 32'h0013469A;
  assign memory[ 2140 ] = 32'h42582100;
  assign memory[ 2141 ] = 32'hE77541A1;
  assign memory[ 2142 ] = 32'h42462700;
  assign memory[ 2143 ] = 32'h2101418F;
  assign memory[ 2144 ] = 32'h468A4249;
  assign memory[ 2145 ] = 32'h42B1E769;
  assign memory[ 2146 ] = 32'hE78ED800;
  assign memory[ 2147 ] = 32'h20002100;
  assign memory[ 2148 ] = 32'h91019000;
  assign memory[ 2149 ] = 32'h29004661;
  assign memory[ 2150 ] = 32'h9800D19E;
  assign memory[ 2151 ] = 32'hE7D39901;
  assign memory[ 2152 ] = 32'h46404662;
  assign memory[ 2153 ] = 32'h46492320;
  assign memory[ 2154 ] = 32'h1A9B4090;
  assign memory[ 2155 ] = 32'h000340D9;
  assign memory[ 2156 ] = 32'h99009100;
  assign memory[ 2157 ] = 32'hE770430B;
  assign memory[ 2158 ] = 32'h23204662;
  assign memory[ 2159 ] = 32'h002A1A9B;
  assign memory[ 2160 ] = 32'h0026409A;
  assign memory[ 2161 ] = 32'h46620013;
  assign memory[ 2162 ] = 32'h431E40D6;
  assign memory[ 2163 ] = 32'h4661E7A9;
  assign memory[ 2164 ] = 32'h27012620;
  assign memory[ 2165 ] = 32'h20001A76;
  assign memory[ 2166 ] = 32'h40F72100;
  assign memory[ 2167 ] = 32'h91019000;
  assign memory[ 2168 ] = 32'hE7729701;
  assign memory[ 2169 ] = 32'h23204662;
  assign memory[ 2170 ] = 32'h40940035;
  assign memory[ 2171 ] = 32'h40DD1A9B;
  assign memory[ 2172 ] = 32'h432B0023;
  assign memory[ 2173 ] = 32'h46C0E79E;
  assign memory[ 2174 ] = 32'h2900B510;
  assign memory[ 2175 ] = 32'hF000D103;
  assign memory[ 2176 ] = 32'h3020F807;
  assign memory[ 2177 ] = 32'h1C08E002;
  assign memory[ 2178 ] = 32'hF802F000;
  assign memory[ 2179 ] = 32'h46C0BD10;
  assign memory[ 2180 ] = 32'h2301211C;
  assign memory[ 2181 ] = 32'h4298041B;
  assign memory[ 2182 ] = 32'h0C00D301;
  assign memory[ 2183 ] = 32'h0A1B3910;
  assign memory[ 2184 ] = 32'hD3014298;
  assign memory[ 2185 ] = 32'h39080A00;
  assign memory[ 2186 ] = 32'h4298091B;
  assign memory[ 2187 ] = 32'h0900D301;
  assign memory[ 2188 ] = 32'hA2023904;
  assign memory[ 2189 ] = 32'h18405C10;
  assign memory[ 2190 ] = 32'h46C04770;
  assign memory[ 2191 ] = 32'h02020304;
  assign memory[ 2192 ] = 32'h01010101;
  assign memory[ 2193 ] = 32'h00000000;
  assign memory[ 2194 ] = 32'h00000000;
  assign memory[ 2195 ] = 32'h0783B570;
  assign memory[ 2196 ] = 32'h1E54D03F;
  assign memory[ 2197 ] = 32'hD03B2A00;
  assign memory[ 2198 ] = 32'h0003B2CE;
  assign memory[ 2199 ] = 32'hE0032503;
  assign memory[ 2200 ] = 32'h2C001E62;
  assign memory[ 2201 ] = 32'h0014D034;
  assign memory[ 2202 ] = 32'h1E5A3301;
  assign memory[ 2203 ] = 32'h422B7016;
  assign memory[ 2204 ] = 32'h2C03D1F6;
  assign memory[ 2205 ] = 32'h25FFD924;
  assign memory[ 2206 ] = 32'h022A400D;
  assign memory[ 2207 ] = 32'h042A4315;
  assign memory[ 2208 ] = 32'h2C0F4315;
  assign memory[ 2209 ] = 32'h0026D911;
  assign memory[ 2210 ] = 32'h09363E10;
  assign memory[ 2211 ] = 32'h01363601;
  assign memory[ 2212 ] = 32'h199B001A;
  assign memory[ 2213 ] = 32'h60556015;
  assign memory[ 2214 ] = 32'h60D56095;
  assign memory[ 2215 ] = 32'h42933210;
  assign memory[ 2216 ] = 32'h220FD1F8;
  assign memory[ 2217 ] = 32'h2C034014;
  assign memory[ 2218 ] = 32'h1F26D90A;
  assign memory[ 2219 ] = 32'h360108B6;
  assign memory[ 2220 ] = 32'h001A00B6;
  assign memory[ 2221 ] = 32'hC220199B;
  assign memory[ 2222 ] = 32'hD1FC4293;
  assign memory[ 2223 ] = 32'h40142203;
  assign memory[ 2224 ] = 32'hD0052C00;
  assign memory[ 2225 ] = 32'h191CB2C9;
  assign memory[ 2226 ] = 32'h33017019;
  assign memory[ 2227 ] = 32'hD1FB429C;
  assign memory[ 2228 ] = 32'h0014BD70;
  assign memory[ 2229 ] = 32'hE7CC0003;
  assign memory[ 2230 ] = 32'h00000676;
  assign memory[ 2231 ] = 32'h00000680;
  assign memory[ 2232 ] = 32'h0000068A;
  assign memory[ 2233 ] = 32'h00000694;
  assign memory[ 2234 ] = 32'h0000069E;
  assign memory[ 2235 ] = 32'h000006A8;
  assign memory[ 2236 ] = 32'h000006B2;
  assign memory[ 2237 ] = 32'h000006BC;
  assign memory[ 2238 ] = 32'h000006C6;
  assign memory[ 2239 ] = 32'h000006D0;
  assign memory[ 2240 ] = 32'h000006DA;
  assign memory[ 2241 ] = 32'h000006E4;
  assign memory[ 2242 ] = 32'h000006EE;
  assign memory[ 2243 ] = 32'h000006F8;
  assign memory[ 2244 ] = 32'h00000702;
  assign memory[ 2245 ] = 32'h0000070C;
  assign memory[ 2246 ] = 32'h40000000;
  assign memory[ 2247 ] = 32'h50000000;
  assign memory[ 2248 ] = 32'h60000000;
  assign memory[ 2249 ] = 32'h00000E9E;
  assign memory[ 2250 ] = 32'h00002A7C;
  assign memory[ 2251 ] = 32'h00000FBA;
  assign memory[ 2252 ] = 32'h00002889;
  assign memory[ 2253 ] = 32'h00001101;
  assign memory[ 2254 ] = 32'h00002A7C;
  assign memory[ 2255 ] = 32'h00001261;
  assign memory[ 2256 ] = 32'h0000248C;
  assign memory[ 2257 ] = 32'h000013DF;
  assign memory[ 2258 ] = 32'h00002281;
  assign memory[ 2259 ] = 32'h0000157C;
  assign memory[ 2260 ] = 32'h0000206F;
  assign memory[ 2261 ] = 32'h0000173A;
  assign memory[ 2262 ] = 32'h00001E56;
  assign memory[ 2263 ] = 32'h0000191B;
  assign memory[ 2264 ] = 32'h00001C35;
  assign memory[ 2265 ] = 32'h00001B24;
  assign memory[ 2266 ] = 32'h00001A0B;
  assign memory[ 2267 ] = 32'h00001D58;
  assign memory[ 2268 ] = 32'h000017D9;
  assign memory[ 2269 ] = 32'h00001FBA;
  assign memory[ 2270 ] = 32'h0000159E;
  assign memory[ 2271 ] = 32'h0000224C;
  assign memory[ 2272 ] = 32'h0000135B;
  assign memory[ 2273 ] = 32'h00002515;
  assign memory[ 2274 ] = 32'h0000110F;
  assign memory[ 2275 ] = 32'h00002817;
  assign memory[ 2276 ] = 32'h00000EBA;
  assign memory[ 2277 ] = 32'h00002B56;
  assign memory[ 2278 ] = 32'h00000C5E;
  assign memory[ 2279 ] = 32'h00002EDB;
  assign memory[ 2280 ] = 32'h000009F6;
  assign memory[ 2281 ] = 32'h000032A6;
  assign memory[ 2282 ] = 32'h00000787;
  assign memory[ 2283 ] = 32'h000036C2;
  assign memory[ 2284 ] = 32'h0000050E;
  assign memory[ 2285 ] = 32'h00003B33;
  assign memory[ 2286 ] = 32'h0000028C;
  assign memory[ 2287 ] = 32'h00004000;
  assign memory[ 2288 ] = 32'h00000000;
  assign memory[ 2289 ] = 32'h0012D687;
  assign memory[ 2290 ] = 32'h00004000;
  assign memory[ 2291 ] = 32'h00000010;
  assign memory[ 2292 ] = 32'h00000666;
  assign memory[ 2293 ] = 32'h0000099A;

// END CUSTOM
 
//Generate the control signals in the address phase
  always_ff @(posedge HCLK, negedge HRESETn)
    if (! HRESETn )
      begin
        read_enable <= '0;
        word_address <= '0;
        byte_select <= '0;
      end
    else if ( HREADY && HSEL && (HTRANS != No_Transfer) )
      begin
        read_enable <= ! HWRITE;
        word_address <= HADDR[MEMWIDTH-1:2];
        byte_select <= generate_byte_select( HSIZE, HADDR[1:0] );
     end
    else
      begin
        read_enable <= '0;
        word_address <= '0;
        byte_select <= '0;
     end

//Act on control signals in the data phase

  // no write since this is a ROM

  //read
  // (output of zero when not enabled for read is not necessary but may help with debugging)
  assign HRDATA[ 7: 0] = ( read_enable && byte_select[0] ) ? memory[word_address][ 7: 0] : '0;
  assign HRDATA[15: 8] = ( read_enable && byte_select[1] ) ? memory[word_address][15: 8] : '0;
  assign HRDATA[23:16] = ( read_enable && byte_select[2] ) ? memory[word_address][23:16] : '0;
  assign HRDATA[31:24] = ( read_enable && byte_select[3] ) ? memory[word_address][31:24] : '0;

//Transfer Response
  assign HREADYOUT = '1; //Single cycle Write & Read. Zero Wait state operations


// decode byte select signals from the size and the lowest two address bits
  function logic [3:0] generate_byte_select( logic [2:0] size, logic [1:0] byte_adress );
    logic byte3, byte2, byte1, byte0;
    byte0 = size[1] || ( byte_adress == 0 );
    byte1 = size[1] || ( size[0] && ( byte_adress == 0 ) ) || ( byte_adress == 1 );
    byte2 = size[1] || ( byte_adress == 2 );
    byte3 = size[1] || ( size[0] && ( byte_adress == 2 ) ) || ( byte_adress == 3 );
    return { byte3, byte2, byte1, byte0 };
  endfunction

endmodule
